-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Nov 17 2024 15:39:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    test : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    test22 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__51921\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51845\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51793\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51764\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51709\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51612\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51600\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51593\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51560\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51548\ : std_logic;
signal \N__51543\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51341\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51230\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51073\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50897\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50894\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50864\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50862\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50843\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50806\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50774\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \N_6_0\ : std_logic;
signal m38 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_120\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_306\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_343_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_344_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.N_43\ : std_logic;
signal \phase_controller_inst1.N_43_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_43_0\ : std_logic;
signal \phase_controller_inst1.running\ : std_logic;
signal \phase_controller_inst1.N_42_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.N_42\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_42_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.start_latched\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.N_38\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.N_38_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.m3_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal s3_phy_c : std_logic;
signal \GB_BUFFER_red_c_g_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.m34_1\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.m10Z0Z_1\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.m3\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.N_1275_i\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.N_139_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.N_34\ : std_logic;
signal \phase_controller_inst2.stoper_hc.m20_nsZ0Z_1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.stoper_hc.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.N_266_0\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_339_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst1.stoper_hc.m19_ns_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_27\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst1.N_175_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_8_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.m12_ns_1\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.N_14_0\ : std_logic;
signal \phase_controller_inst1.N_13_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.m21\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.time_passed_er_RNI23UO1\ : std_logic;
signal s1_phy_c : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_45_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \S1_RNI9RLH\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_286\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_339_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_8_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal test22_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_340_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_287_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_45\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_46\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_46_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_46_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_342_i\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.N_265_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.N_47\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.mZ0Z16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.m28_ns_1\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \GNDG0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_5\ : std_logic;
signal test_c : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.start_latched\ : std_logic;
signal \phase_controller_inst2.running\ : std_logic;
signal \phase_controller_inst2.N_39\ : std_logic;
signal \phase_controller_inst2.stoper_tr.N_39_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_289\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_290\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_341_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal clock_output_0 : std_logic;
signal red_c_g : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal test_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal test22_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    test <= test_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    test22 <= test22_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__37148\&\N__37188\&\N__37230\&\N__37274\&\N__37317\&\N__36822\&\N__36870\&\N__36906\&\N__36938\&\N__36984\&\N__37022\&\N__37059\&\N__36494\&\N__36531\&\N__36579\&\N__36612\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__49818\&'0'&\N__49817\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21601\&\N__21594\&\N__21599\&\N__21593\&\N__21600\&\N__21592\&\N__21602\&\N__21589\&\N__21595\&\N__21588\&\N__21596\&\N__21590\&\N__21597\&\N__21591\&\N__21598\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__49871\&\N__49868\&'0'&'0'&'0'&\N__49866\&\N__49870\&\N__49867\&\N__49869\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21562\&\N__21565\&\N__21563\&\N__21566\&\N__21564\&\N__19483\&\N__19498\&\N__19463\&\N__19441\&\N__19425\&\N__20517\&\N__20542\&\N__19272\&\N__19287\&\N__19302\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__49796\&\N__49793\&'0'&'0'&'0'&\N__49791\&\N__49795\&\N__49792\&\N__49794\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__36644\&\N__36680\&\N__36726\&\N__36768\&\N__36240\&\N__36282\&\N__38229\&\N__36321\&\N__36363\&\N__36395\&\N__50967\&\N__36450\&\N__35970\&\N__36015\&\N__30695\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__49660\&'0'&\N__49659\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__25797\,
            RESETB => \N__31242\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__49826\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__49816\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__49872\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__49865\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__49797\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__49790\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__49825\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__49658\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__51919\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51921\,
            DIN => \N__51920\,
            DOUT => \N__51919\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51921\,
            PADOUT => \N__51920\,
            PADIN => \N__51919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51910\,
            DIN => \N__51909\,
            DOUT => \N__51908\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51910\,
            PADOUT => \N__51909\,
            PADIN => \N__51908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__47493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51901\,
            DIN => \N__51900\,
            DOUT => \N__51899\,
            PACKAGEPIN => test_wire
        );

    \test_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51901\,
            PADOUT => \N__51900\,
            PADIN => \N__51899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43701\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51892\,
            DIN => \N__51891\,
            DOUT => \N__51890\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51892\,
            PADOUT => \N__51891\,
            PADIN => \N__51890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51883\,
            DIN => \N__51882\,
            DOUT => \N__51881\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51883\,
            PADOUT => \N__51882\,
            PADIN => \N__51881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51874\,
            DIN => \N__51873\,
            DOUT => \N__51872\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51874\,
            PADOUT => \N__51873\,
            PADIN => \N__51872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21750\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51865\,
            DIN => \N__51864\,
            DOUT => \N__51863\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51865\,
            PADOUT => \N__51864\,
            PADIN => \N__51863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51856\,
            DIN => \N__51855\,
            DOUT => \N__51854\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51856\,
            PADOUT => \N__51855\,
            PADIN => \N__51854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37086\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test22_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51847\,
            DIN => \N__51846\,
            DOUT => \N__51845\,
            PACKAGEPIN => test22_wire
        );

    \test22_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51847\,
            PADOUT => \N__51846\,
            PADIN => \N__51845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38745\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51838\,
            DIN => \N__51837\,
            DOUT => \N__51836\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51838\,
            PADOUT => \N__51837\,
            PADIN => \N__51836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51829\,
            DIN => \N__51828\,
            DOUT => \N__51827\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51829\,
            PADOUT => \N__51828\,
            PADIN => \N__51827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51820\,
            DIN => \N__51819\,
            DOUT => \N__51818\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51820\,
            PADOUT => \N__51819\,
            PADIN => \N__51818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51811\,
            DIN => \N__51810\,
            DOUT => \N__51809\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51811\,
            PADOUT => \N__51810\,
            PADIN => \N__51809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51802\,
            DIN => \N__51801\,
            DOUT => \N__51800\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51802\,
            PADOUT => \N__51801\,
            PADIN => \N__51800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31257\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51793\,
            DIN => \N__51792\,
            DOUT => \N__51791\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51793\,
            PADOUT => \N__51792\,
            PADIN => \N__51791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51784\,
            DIN => \N__51783\,
            DOUT => \N__51782\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__51784\,
            PADOUT => \N__51783\,
            PADIN => \N__51782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12456\ : InMux
    port map (
            O => \N__51765\,
            I => \N__51759\
        );

    \I__12455\ : InMux
    port map (
            O => \N__51764\,
            I => \N__51756\
        );

    \I__12454\ : InMux
    port map (
            O => \N__51763\,
            I => \N__51753\
        );

    \I__12453\ : InMux
    port map (
            O => \N__51762\,
            I => \N__51750\
        );

    \I__12452\ : LocalMux
    port map (
            O => \N__51759\,
            I => \N__51747\
        );

    \I__12451\ : LocalMux
    port map (
            O => \N__51756\,
            I => \N__51744\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__51753\,
            I => \N__51741\
        );

    \I__12449\ : LocalMux
    port map (
            O => \N__51750\,
            I => \N__51738\
        );

    \I__12448\ : Span4Mux_h
    port map (
            O => \N__51747\,
            I => \N__51735\
        );

    \I__12447\ : Span4Mux_h
    port map (
            O => \N__51744\,
            I => \N__51730\
        );

    \I__12446\ : Span4Mux_h
    port map (
            O => \N__51741\,
            I => \N__51730\
        );

    \I__12445\ : Odrv4
    port map (
            O => \N__51738\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__12444\ : Odrv4
    port map (
            O => \N__51735\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__12443\ : Odrv4
    port map (
            O => \N__51730\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__12442\ : InMux
    port map (
            O => \N__51723\,
            I => \N__51720\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__51720\,
            I => \N__51717\
        );

    \I__12440\ : Span4Mux_v
    port map (
            O => \N__51717\,
            I => \N__51712\
        );

    \I__12439\ : InMux
    port map (
            O => \N__51716\,
            I => \N__51709\
        );

    \I__12438\ : InMux
    port map (
            O => \N__51715\,
            I => \N__51706\
        );

    \I__12437\ : Span4Mux_h
    port map (
            O => \N__51712\,
            I => \N__51701\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__51709\,
            I => \N__51701\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__51706\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__12434\ : Odrv4
    port map (
            O => \N__51701\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__12433\ : InMux
    port map (
            O => \N__51696\,
            I => \N__51690\
        );

    \I__12432\ : InMux
    port map (
            O => \N__51695\,
            I => \N__51687\
        );

    \I__12431\ : InMux
    port map (
            O => \N__51694\,
            I => \N__51684\
        );

    \I__12430\ : InMux
    port map (
            O => \N__51693\,
            I => \N__51681\
        );

    \I__12429\ : LocalMux
    port map (
            O => \N__51690\,
            I => \N__51678\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__51687\,
            I => \N__51675\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__51684\,
            I => \N__51672\
        );

    \I__12426\ : LocalMux
    port map (
            O => \N__51681\,
            I => \N__51669\
        );

    \I__12425\ : Span4Mux_v
    port map (
            O => \N__51678\,
            I => \N__51664\
        );

    \I__12424\ : Span4Mux_v
    port map (
            O => \N__51675\,
            I => \N__51664\
        );

    \I__12423\ : Span4Mux_h
    port map (
            O => \N__51672\,
            I => \N__51661\
        );

    \I__12422\ : Odrv12
    port map (
            O => \N__51669\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__12421\ : Odrv4
    port map (
            O => \N__51664\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__12420\ : Odrv4
    port map (
            O => \N__51661\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__12419\ : InMux
    port map (
            O => \N__51654\,
            I => \N__51650\
        );

    \I__12418\ : InMux
    port map (
            O => \N__51653\,
            I => \N__51647\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__51650\,
            I => \N__51643\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__51647\,
            I => \N__51640\
        );

    \I__12415\ : InMux
    port map (
            O => \N__51646\,
            I => \N__51637\
        );

    \I__12414\ : Span4Mux_h
    port map (
            O => \N__51643\,
            I => \N__51634\
        );

    \I__12413\ : Span4Mux_v
    port map (
            O => \N__51640\,
            I => \N__51631\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__51637\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12411\ : Odrv4
    port map (
            O => \N__51634\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12410\ : Odrv4
    port map (
            O => \N__51631\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12409\ : CascadeMux
    port map (
            O => \N__51624\,
            I => \N__51613\
        );

    \I__12408\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51605\
        );

    \I__12407\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51605\
        );

    \I__12406\ : InMux
    port map (
            O => \N__51621\,
            I => \N__51605\
        );

    \I__12405\ : InMux
    port map (
            O => \N__51620\,
            I => \N__51597\
        );

    \I__12404\ : InMux
    port map (
            O => \N__51619\,
            I => \N__51589\
        );

    \I__12403\ : InMux
    port map (
            O => \N__51618\,
            I => \N__51582\
        );

    \I__12402\ : InMux
    port map (
            O => \N__51617\,
            I => \N__51582\
        );

    \I__12401\ : InMux
    port map (
            O => \N__51616\,
            I => \N__51582\
        );

    \I__12400\ : InMux
    port map (
            O => \N__51613\,
            I => \N__51574\
        );

    \I__12399\ : InMux
    port map (
            O => \N__51612\,
            I => \N__51574\
        );

    \I__12398\ : LocalMux
    port map (
            O => \N__51605\,
            I => \N__51571\
        );

    \I__12397\ : InMux
    port map (
            O => \N__51604\,
            I => \N__51560\
        );

    \I__12396\ : InMux
    port map (
            O => \N__51603\,
            I => \N__51560\
        );

    \I__12395\ : InMux
    port map (
            O => \N__51602\,
            I => \N__51560\
        );

    \I__12394\ : InMux
    port map (
            O => \N__51601\,
            I => \N__51560\
        );

    \I__12393\ : InMux
    port map (
            O => \N__51600\,
            I => \N__51560\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__51597\,
            I => \N__51548\
        );

    \I__12391\ : InMux
    port map (
            O => \N__51596\,
            I => \N__51543\
        );

    \I__12390\ : InMux
    port map (
            O => \N__51595\,
            I => \N__51543\
        );

    \I__12389\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51536\
        );

    \I__12388\ : InMux
    port map (
            O => \N__51593\,
            I => \N__51536\
        );

    \I__12387\ : InMux
    port map (
            O => \N__51592\,
            I => \N__51536\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__51589\,
            I => \N__51531\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__51582\,
            I => \N__51531\
        );

    \I__12384\ : InMux
    port map (
            O => \N__51581\,
            I => \N__51526\
        );

    \I__12383\ : InMux
    port map (
            O => \N__51580\,
            I => \N__51526\
        );

    \I__12382\ : CascadeMux
    port map (
            O => \N__51579\,
            I => \N__51523\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__51574\,
            I => \N__51508\
        );

    \I__12380\ : Span4Mux_v
    port map (
            O => \N__51571\,
            I => \N__51508\
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__51560\,
            I => \N__51508\
        );

    \I__12378\ : InMux
    port map (
            O => \N__51559\,
            I => \N__51505\
        );

    \I__12377\ : InMux
    port map (
            O => \N__51558\,
            I => \N__51494\
        );

    \I__12376\ : InMux
    port map (
            O => \N__51557\,
            I => \N__51494\
        );

    \I__12375\ : InMux
    port map (
            O => \N__51556\,
            I => \N__51494\
        );

    \I__12374\ : InMux
    port map (
            O => \N__51555\,
            I => \N__51491\
        );

    \I__12373\ : InMux
    port map (
            O => \N__51554\,
            I => \N__51488\
        );

    \I__12372\ : InMux
    port map (
            O => \N__51553\,
            I => \N__51483\
        );

    \I__12371\ : InMux
    port map (
            O => \N__51552\,
            I => \N__51483\
        );

    \I__12370\ : InMux
    port map (
            O => \N__51551\,
            I => \N__51480\
        );

    \I__12369\ : Span4Mux_v
    port map (
            O => \N__51548\,
            I => \N__51469\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__51543\,
            I => \N__51469\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__51536\,
            I => \N__51469\
        );

    \I__12366\ : Span4Mux_v
    port map (
            O => \N__51531\,
            I => \N__51469\
        );

    \I__12365\ : LocalMux
    port map (
            O => \N__51526\,
            I => \N__51469\
        );

    \I__12364\ : InMux
    port map (
            O => \N__51523\,
            I => \N__51464\
        );

    \I__12363\ : InMux
    port map (
            O => \N__51522\,
            I => \N__51464\
        );

    \I__12362\ : InMux
    port map (
            O => \N__51521\,
            I => \N__51461\
        );

    \I__12361\ : CascadeMux
    port map (
            O => \N__51520\,
            I => \N__51457\
        );

    \I__12360\ : InMux
    port map (
            O => \N__51519\,
            I => \N__51450\
        );

    \I__12359\ : InMux
    port map (
            O => \N__51518\,
            I => \N__51450\
        );

    \I__12358\ : InMux
    port map (
            O => \N__51517\,
            I => \N__51450\
        );

    \I__12357\ : CascadeMux
    port map (
            O => \N__51516\,
            I => \N__51447\
        );

    \I__12356\ : InMux
    port map (
            O => \N__51515\,
            I => \N__51427\
        );

    \I__12355\ : Span4Mux_v
    port map (
            O => \N__51508\,
            I => \N__51422\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__51505\,
            I => \N__51422\
        );

    \I__12353\ : InMux
    port map (
            O => \N__51504\,
            I => \N__51419\
        );

    \I__12352\ : InMux
    port map (
            O => \N__51503\,
            I => \N__51416\
        );

    \I__12351\ : InMux
    port map (
            O => \N__51502\,
            I => \N__51410\
        );

    \I__12350\ : InMux
    port map (
            O => \N__51501\,
            I => \N__51410\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__51494\,
            I => \N__51395\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__51491\,
            I => \N__51395\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__51488\,
            I => \N__51395\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__51483\,
            I => \N__51395\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__51480\,
            I => \N__51395\
        );

    \I__12344\ : Span4Mux_v
    port map (
            O => \N__51469\,
            I => \N__51395\
        );

    \I__12343\ : LocalMux
    port map (
            O => \N__51464\,
            I => \N__51395\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__51461\,
            I => \N__51392\
        );

    \I__12341\ : CascadeMux
    port map (
            O => \N__51460\,
            I => \N__51383\
        );

    \I__12340\ : InMux
    port map (
            O => \N__51457\,
            I => \N__51380\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__51450\,
            I => \N__51377\
        );

    \I__12338\ : InMux
    port map (
            O => \N__51447\,
            I => \N__51374\
        );

    \I__12337\ : InMux
    port map (
            O => \N__51446\,
            I => \N__51369\
        );

    \I__12336\ : InMux
    port map (
            O => \N__51445\,
            I => \N__51369\
        );

    \I__12335\ : InMux
    port map (
            O => \N__51444\,
            I => \N__51362\
        );

    \I__12334\ : InMux
    port map (
            O => \N__51443\,
            I => \N__51362\
        );

    \I__12333\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51362\
        );

    \I__12332\ : InMux
    port map (
            O => \N__51441\,
            I => \N__51351\
        );

    \I__12331\ : InMux
    port map (
            O => \N__51440\,
            I => \N__51351\
        );

    \I__12330\ : InMux
    port map (
            O => \N__51439\,
            I => \N__51351\
        );

    \I__12329\ : InMux
    port map (
            O => \N__51438\,
            I => \N__51351\
        );

    \I__12328\ : InMux
    port map (
            O => \N__51437\,
            I => \N__51351\
        );

    \I__12327\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51346\
        );

    \I__12326\ : InMux
    port map (
            O => \N__51435\,
            I => \N__51346\
        );

    \I__12325\ : InMux
    port map (
            O => \N__51434\,
            I => \N__51341\
        );

    \I__12324\ : InMux
    port map (
            O => \N__51433\,
            I => \N__51341\
        );

    \I__12323\ : InMux
    port map (
            O => \N__51432\,
            I => \N__51336\
        );

    \I__12322\ : InMux
    port map (
            O => \N__51431\,
            I => \N__51336\
        );

    \I__12321\ : InMux
    port map (
            O => \N__51430\,
            I => \N__51333\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__51427\,
            I => \N__51326\
        );

    \I__12319\ : Span4Mux_h
    port map (
            O => \N__51422\,
            I => \N__51326\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__51419\,
            I => \N__51326\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__51416\,
            I => \N__51323\
        );

    \I__12316\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51310\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__51410\,
            I => \N__51307\
        );

    \I__12314\ : Span4Mux_v
    port map (
            O => \N__51395\,
            I => \N__51302\
        );

    \I__12313\ : Span4Mux_v
    port map (
            O => \N__51392\,
            I => \N__51302\
        );

    \I__12312\ : InMux
    port map (
            O => \N__51391\,
            I => \N__51289\
        );

    \I__12311\ : InMux
    port map (
            O => \N__51390\,
            I => \N__51289\
        );

    \I__12310\ : InMux
    port map (
            O => \N__51389\,
            I => \N__51289\
        );

    \I__12309\ : InMux
    port map (
            O => \N__51388\,
            I => \N__51289\
        );

    \I__12308\ : InMux
    port map (
            O => \N__51387\,
            I => \N__51275\
        );

    \I__12307\ : InMux
    port map (
            O => \N__51386\,
            I => \N__51275\
        );

    \I__12306\ : InMux
    port map (
            O => \N__51383\,
            I => \N__51272\
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__51380\,
            I => \N__51269\
        );

    \I__12304\ : Span4Mux_h
    port map (
            O => \N__51377\,
            I => \N__51264\
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__51374\,
            I => \N__51264\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__51369\,
            I => \N__51261\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__51362\,
            I => \N__51254\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__51351\,
            I => \N__51254\
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__51346\,
            I => \N__51254\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__51341\,
            I => \N__51251\
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__51336\,
            I => \N__51242\
        );

    \I__12296\ : LocalMux
    port map (
            O => \N__51333\,
            I => \N__51242\
        );

    \I__12295\ : Span4Mux_v
    port map (
            O => \N__51326\,
            I => \N__51242\
        );

    \I__12294\ : Span4Mux_v
    port map (
            O => \N__51323\,
            I => \N__51242\
        );

    \I__12293\ : InMux
    port map (
            O => \N__51322\,
            I => \N__51233\
        );

    \I__12292\ : InMux
    port map (
            O => \N__51321\,
            I => \N__51233\
        );

    \I__12291\ : InMux
    port map (
            O => \N__51320\,
            I => \N__51233\
        );

    \I__12290\ : InMux
    port map (
            O => \N__51319\,
            I => \N__51233\
        );

    \I__12289\ : InMux
    port map (
            O => \N__51318\,
            I => \N__51230\
        );

    \I__12288\ : InMux
    port map (
            O => \N__51317\,
            I => \N__51227\
        );

    \I__12287\ : InMux
    port map (
            O => \N__51316\,
            I => \N__51218\
        );

    \I__12286\ : InMux
    port map (
            O => \N__51315\,
            I => \N__51218\
        );

    \I__12285\ : InMux
    port map (
            O => \N__51314\,
            I => \N__51218\
        );

    \I__12284\ : InMux
    port map (
            O => \N__51313\,
            I => \N__51218\
        );

    \I__12283\ : LocalMux
    port map (
            O => \N__51310\,
            I => \N__51211\
        );

    \I__12282\ : Span4Mux_v
    port map (
            O => \N__51307\,
            I => \N__51211\
        );

    \I__12281\ : Span4Mux_h
    port map (
            O => \N__51302\,
            I => \N__51211\
        );

    \I__12280\ : InMux
    port map (
            O => \N__51301\,
            I => \N__51206\
        );

    \I__12279\ : InMux
    port map (
            O => \N__51300\,
            I => \N__51206\
        );

    \I__12278\ : InMux
    port map (
            O => \N__51299\,
            I => \N__51203\
        );

    \I__12277\ : InMux
    port map (
            O => \N__51298\,
            I => \N__51200\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__51289\,
            I => \N__51197\
        );

    \I__12275\ : InMux
    port map (
            O => \N__51288\,
            I => \N__51190\
        );

    \I__12274\ : InMux
    port map (
            O => \N__51287\,
            I => \N__51190\
        );

    \I__12273\ : InMux
    port map (
            O => \N__51286\,
            I => \N__51190\
        );

    \I__12272\ : InMux
    port map (
            O => \N__51285\,
            I => \N__51183\
        );

    \I__12271\ : InMux
    port map (
            O => \N__51284\,
            I => \N__51183\
        );

    \I__12270\ : InMux
    port map (
            O => \N__51283\,
            I => \N__51183\
        );

    \I__12269\ : InMux
    port map (
            O => \N__51282\,
            I => \N__51176\
        );

    \I__12268\ : InMux
    port map (
            O => \N__51281\,
            I => \N__51176\
        );

    \I__12267\ : InMux
    port map (
            O => \N__51280\,
            I => \N__51176\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__51275\,
            I => \N__51159\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__51272\,
            I => \N__51159\
        );

    \I__12264\ : Span4Mux_v
    port map (
            O => \N__51269\,
            I => \N__51159\
        );

    \I__12263\ : Span4Mux_v
    port map (
            O => \N__51264\,
            I => \N__51159\
        );

    \I__12262\ : Span4Mux_v
    port map (
            O => \N__51261\,
            I => \N__51159\
        );

    \I__12261\ : Span4Mux_v
    port map (
            O => \N__51254\,
            I => \N__51159\
        );

    \I__12260\ : Span4Mux_h
    port map (
            O => \N__51251\,
            I => \N__51159\
        );

    \I__12259\ : Span4Mux_h
    port map (
            O => \N__51242\,
            I => \N__51159\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__51233\,
            I => \N__51148\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__51230\,
            I => \N__51148\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__51227\,
            I => \N__51148\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__51218\,
            I => \N__51148\
        );

    \I__12254\ : Span4Mux_v
    port map (
            O => \N__51211\,
            I => \N__51148\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__51206\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__51203\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__51200\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12250\ : Odrv4
    port map (
            O => \N__51197\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__51190\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__51183\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__51176\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12246\ : Odrv4
    port map (
            O => \N__51159\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12245\ : Odrv4
    port map (
            O => \N__51148\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__12244\ : InMux
    port map (
            O => \N__51129\,
            I => \N__51124\
        );

    \I__12243\ : InMux
    port map (
            O => \N__51128\,
            I => \N__51120\
        );

    \I__12242\ : InMux
    port map (
            O => \N__51127\,
            I => \N__51117\
        );

    \I__12241\ : LocalMux
    port map (
            O => \N__51124\,
            I => \N__51114\
        );

    \I__12240\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51111\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__51120\,
            I => \N__51108\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__51117\,
            I => \N__51103\
        );

    \I__12237\ : Span4Mux_v
    port map (
            O => \N__51114\,
            I => \N__51103\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__51111\,
            I => \N__51100\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__51108\,
            I => \N__51097\
        );

    \I__12234\ : Span4Mux_h
    port map (
            O => \N__51103\,
            I => \N__51092\
        );

    \I__12233\ : Span4Mux_h
    port map (
            O => \N__51100\,
            I => \N__51092\
        );

    \I__12232\ : Odrv4
    port map (
            O => \N__51097\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__12231\ : Odrv4
    port map (
            O => \N__51092\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__12230\ : InMux
    port map (
            O => \N__51087\,
            I => \N__51083\
        );

    \I__12229\ : InMux
    port map (
            O => \N__51086\,
            I => \N__51079\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__51083\,
            I => \N__51076\
        );

    \I__12227\ : InMux
    port map (
            O => \N__51082\,
            I => \N__51073\
        );

    \I__12226\ : LocalMux
    port map (
            O => \N__51079\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__12225\ : Odrv4
    port map (
            O => \N__51076\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__51073\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__12223\ : InMux
    port map (
            O => \N__51066\,
            I => \N__51062\
        );

    \I__12222\ : InMux
    port map (
            O => \N__51065\,
            I => \N__51059\
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__51062\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__51059\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__12219\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51051\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__51051\,
            I => \N__51047\
        );

    \I__12217\ : InMux
    port map (
            O => \N__51050\,
            I => \N__51044\
        );

    \I__12216\ : Span4Mux_h
    port map (
            O => \N__51047\,
            I => \N__51038\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__51044\,
            I => \N__51038\
        );

    \I__12214\ : InMux
    port map (
            O => \N__51043\,
            I => \N__51035\
        );

    \I__12213\ : Span4Mux_h
    port map (
            O => \N__51038\,
            I => \N__51032\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__51035\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__12211\ : Odrv4
    port map (
            O => \N__51032\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__12210\ : CascadeMux
    port map (
            O => \N__51027\,
            I => \N__51023\
        );

    \I__12209\ : CascadeMux
    port map (
            O => \N__51026\,
            I => \N__51020\
        );

    \I__12208\ : InMux
    port map (
            O => \N__51023\,
            I => \N__51017\
        );

    \I__12207\ : InMux
    port map (
            O => \N__51020\,
            I => \N__51014\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__51017\,
            I => \N__51008\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__51014\,
            I => \N__51008\
        );

    \I__12204\ : InMux
    port map (
            O => \N__51013\,
            I => \N__51005\
        );

    \I__12203\ : Span4Mux_v
    port map (
            O => \N__51008\,
            I => \N__51002\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__51005\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__12201\ : Odrv4
    port map (
            O => \N__51002\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__12200\ : InMux
    port map (
            O => \N__50997\,
            I => \N__50993\
        );

    \I__12199\ : InMux
    port map (
            O => \N__50996\,
            I => \N__50990\
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__50993\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__12197\ : LocalMux
    port map (
            O => \N__50990\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__12196\ : CascadeMux
    port map (
            O => \N__50985\,
            I => \N__50982\
        );

    \I__12195\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50979\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__50979\,
            I => \N__50976\
        );

    \I__12193\ : Span4Mux_h
    port map (
            O => \N__50976\,
            I => \N__50973\
        );

    \I__12192\ : Span4Mux_v
    port map (
            O => \N__50973\,
            I => \N__50970\
        );

    \I__12191\ : Odrv4
    port map (
            O => \N__50970\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__12190\ : InMux
    port map (
            O => \N__50967\,
            I => \N__50963\
        );

    \I__12189\ : InMux
    port map (
            O => \N__50966\,
            I => \N__50960\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__50963\,
            I => \N__50957\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__50960\,
            I => \N__50954\
        );

    \I__12186\ : Span4Mux_v
    port map (
            O => \N__50957\,
            I => \N__50951\
        );

    \I__12185\ : Span4Mux_v
    port map (
            O => \N__50954\,
            I => \N__50946\
        );

    \I__12184\ : Span4Mux_v
    port map (
            O => \N__50951\,
            I => \N__50946\
        );

    \I__12183\ : Sp12to4
    port map (
            O => \N__50946\,
            I => \N__50943\
        );

    \I__12182\ : Odrv12
    port map (
            O => \N__50943\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__12181\ : InMux
    port map (
            O => \N__50940\,
            I => \N__50937\
        );

    \I__12180\ : LocalMux
    port map (
            O => \N__50937\,
            I => \N__50934\
        );

    \I__12179\ : Span4Mux_h
    port map (
            O => \N__50934\,
            I => \N__50931\
        );

    \I__12178\ : Span4Mux_h
    port map (
            O => \N__50931\,
            I => \N__50928\
        );

    \I__12177\ : Span4Mux_h
    port map (
            O => \N__50928\,
            I => \N__50925\
        );

    \I__12176\ : Span4Mux_h
    port map (
            O => \N__50925\,
            I => \N__50922\
        );

    \I__12175\ : Odrv4
    port map (
            O => \N__50922\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__12174\ : InMux
    port map (
            O => \N__50919\,
            I => \N__50916\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__50916\,
            I => \N__50753\
        );

    \I__12172\ : ClkMux
    port map (
            O => \N__50915\,
            I => \N__50421\
        );

    \I__12171\ : ClkMux
    port map (
            O => \N__50914\,
            I => \N__50421\
        );

    \I__12170\ : ClkMux
    port map (
            O => \N__50913\,
            I => \N__50421\
        );

    \I__12169\ : ClkMux
    port map (
            O => \N__50912\,
            I => \N__50421\
        );

    \I__12168\ : ClkMux
    port map (
            O => \N__50911\,
            I => \N__50421\
        );

    \I__12167\ : ClkMux
    port map (
            O => \N__50910\,
            I => \N__50421\
        );

    \I__12166\ : ClkMux
    port map (
            O => \N__50909\,
            I => \N__50421\
        );

    \I__12165\ : ClkMux
    port map (
            O => \N__50908\,
            I => \N__50421\
        );

    \I__12164\ : ClkMux
    port map (
            O => \N__50907\,
            I => \N__50421\
        );

    \I__12163\ : ClkMux
    port map (
            O => \N__50906\,
            I => \N__50421\
        );

    \I__12162\ : ClkMux
    port map (
            O => \N__50905\,
            I => \N__50421\
        );

    \I__12161\ : ClkMux
    port map (
            O => \N__50904\,
            I => \N__50421\
        );

    \I__12160\ : ClkMux
    port map (
            O => \N__50903\,
            I => \N__50421\
        );

    \I__12159\ : ClkMux
    port map (
            O => \N__50902\,
            I => \N__50421\
        );

    \I__12158\ : ClkMux
    port map (
            O => \N__50901\,
            I => \N__50421\
        );

    \I__12157\ : ClkMux
    port map (
            O => \N__50900\,
            I => \N__50421\
        );

    \I__12156\ : ClkMux
    port map (
            O => \N__50899\,
            I => \N__50421\
        );

    \I__12155\ : ClkMux
    port map (
            O => \N__50898\,
            I => \N__50421\
        );

    \I__12154\ : ClkMux
    port map (
            O => \N__50897\,
            I => \N__50421\
        );

    \I__12153\ : ClkMux
    port map (
            O => \N__50896\,
            I => \N__50421\
        );

    \I__12152\ : ClkMux
    port map (
            O => \N__50895\,
            I => \N__50421\
        );

    \I__12151\ : ClkMux
    port map (
            O => \N__50894\,
            I => \N__50421\
        );

    \I__12150\ : ClkMux
    port map (
            O => \N__50893\,
            I => \N__50421\
        );

    \I__12149\ : ClkMux
    port map (
            O => \N__50892\,
            I => \N__50421\
        );

    \I__12148\ : ClkMux
    port map (
            O => \N__50891\,
            I => \N__50421\
        );

    \I__12147\ : ClkMux
    port map (
            O => \N__50890\,
            I => \N__50421\
        );

    \I__12146\ : ClkMux
    port map (
            O => \N__50889\,
            I => \N__50421\
        );

    \I__12145\ : ClkMux
    port map (
            O => \N__50888\,
            I => \N__50421\
        );

    \I__12144\ : ClkMux
    port map (
            O => \N__50887\,
            I => \N__50421\
        );

    \I__12143\ : ClkMux
    port map (
            O => \N__50886\,
            I => \N__50421\
        );

    \I__12142\ : ClkMux
    port map (
            O => \N__50885\,
            I => \N__50421\
        );

    \I__12141\ : ClkMux
    port map (
            O => \N__50884\,
            I => \N__50421\
        );

    \I__12140\ : ClkMux
    port map (
            O => \N__50883\,
            I => \N__50421\
        );

    \I__12139\ : ClkMux
    port map (
            O => \N__50882\,
            I => \N__50421\
        );

    \I__12138\ : ClkMux
    port map (
            O => \N__50881\,
            I => \N__50421\
        );

    \I__12137\ : ClkMux
    port map (
            O => \N__50880\,
            I => \N__50421\
        );

    \I__12136\ : ClkMux
    port map (
            O => \N__50879\,
            I => \N__50421\
        );

    \I__12135\ : ClkMux
    port map (
            O => \N__50878\,
            I => \N__50421\
        );

    \I__12134\ : ClkMux
    port map (
            O => \N__50877\,
            I => \N__50421\
        );

    \I__12133\ : ClkMux
    port map (
            O => \N__50876\,
            I => \N__50421\
        );

    \I__12132\ : ClkMux
    port map (
            O => \N__50875\,
            I => \N__50421\
        );

    \I__12131\ : ClkMux
    port map (
            O => \N__50874\,
            I => \N__50421\
        );

    \I__12130\ : ClkMux
    port map (
            O => \N__50873\,
            I => \N__50421\
        );

    \I__12129\ : ClkMux
    port map (
            O => \N__50872\,
            I => \N__50421\
        );

    \I__12128\ : ClkMux
    port map (
            O => \N__50871\,
            I => \N__50421\
        );

    \I__12127\ : ClkMux
    port map (
            O => \N__50870\,
            I => \N__50421\
        );

    \I__12126\ : ClkMux
    port map (
            O => \N__50869\,
            I => \N__50421\
        );

    \I__12125\ : ClkMux
    port map (
            O => \N__50868\,
            I => \N__50421\
        );

    \I__12124\ : ClkMux
    port map (
            O => \N__50867\,
            I => \N__50421\
        );

    \I__12123\ : ClkMux
    port map (
            O => \N__50866\,
            I => \N__50421\
        );

    \I__12122\ : ClkMux
    port map (
            O => \N__50865\,
            I => \N__50421\
        );

    \I__12121\ : ClkMux
    port map (
            O => \N__50864\,
            I => \N__50421\
        );

    \I__12120\ : ClkMux
    port map (
            O => \N__50863\,
            I => \N__50421\
        );

    \I__12119\ : ClkMux
    port map (
            O => \N__50862\,
            I => \N__50421\
        );

    \I__12118\ : ClkMux
    port map (
            O => \N__50861\,
            I => \N__50421\
        );

    \I__12117\ : ClkMux
    port map (
            O => \N__50860\,
            I => \N__50421\
        );

    \I__12116\ : ClkMux
    port map (
            O => \N__50859\,
            I => \N__50421\
        );

    \I__12115\ : ClkMux
    port map (
            O => \N__50858\,
            I => \N__50421\
        );

    \I__12114\ : ClkMux
    port map (
            O => \N__50857\,
            I => \N__50421\
        );

    \I__12113\ : ClkMux
    port map (
            O => \N__50856\,
            I => \N__50421\
        );

    \I__12112\ : ClkMux
    port map (
            O => \N__50855\,
            I => \N__50421\
        );

    \I__12111\ : ClkMux
    port map (
            O => \N__50854\,
            I => \N__50421\
        );

    \I__12110\ : ClkMux
    port map (
            O => \N__50853\,
            I => \N__50421\
        );

    \I__12109\ : ClkMux
    port map (
            O => \N__50852\,
            I => \N__50421\
        );

    \I__12108\ : ClkMux
    port map (
            O => \N__50851\,
            I => \N__50421\
        );

    \I__12107\ : ClkMux
    port map (
            O => \N__50850\,
            I => \N__50421\
        );

    \I__12106\ : ClkMux
    port map (
            O => \N__50849\,
            I => \N__50421\
        );

    \I__12105\ : ClkMux
    port map (
            O => \N__50848\,
            I => \N__50421\
        );

    \I__12104\ : ClkMux
    port map (
            O => \N__50847\,
            I => \N__50421\
        );

    \I__12103\ : ClkMux
    port map (
            O => \N__50846\,
            I => \N__50421\
        );

    \I__12102\ : ClkMux
    port map (
            O => \N__50845\,
            I => \N__50421\
        );

    \I__12101\ : ClkMux
    port map (
            O => \N__50844\,
            I => \N__50421\
        );

    \I__12100\ : ClkMux
    port map (
            O => \N__50843\,
            I => \N__50421\
        );

    \I__12099\ : ClkMux
    port map (
            O => \N__50842\,
            I => \N__50421\
        );

    \I__12098\ : ClkMux
    port map (
            O => \N__50841\,
            I => \N__50421\
        );

    \I__12097\ : ClkMux
    port map (
            O => \N__50840\,
            I => \N__50421\
        );

    \I__12096\ : ClkMux
    port map (
            O => \N__50839\,
            I => \N__50421\
        );

    \I__12095\ : ClkMux
    port map (
            O => \N__50838\,
            I => \N__50421\
        );

    \I__12094\ : ClkMux
    port map (
            O => \N__50837\,
            I => \N__50421\
        );

    \I__12093\ : ClkMux
    port map (
            O => \N__50836\,
            I => \N__50421\
        );

    \I__12092\ : ClkMux
    port map (
            O => \N__50835\,
            I => \N__50421\
        );

    \I__12091\ : ClkMux
    port map (
            O => \N__50834\,
            I => \N__50421\
        );

    \I__12090\ : ClkMux
    port map (
            O => \N__50833\,
            I => \N__50421\
        );

    \I__12089\ : ClkMux
    port map (
            O => \N__50832\,
            I => \N__50421\
        );

    \I__12088\ : ClkMux
    port map (
            O => \N__50831\,
            I => \N__50421\
        );

    \I__12087\ : ClkMux
    port map (
            O => \N__50830\,
            I => \N__50421\
        );

    \I__12086\ : ClkMux
    port map (
            O => \N__50829\,
            I => \N__50421\
        );

    \I__12085\ : ClkMux
    port map (
            O => \N__50828\,
            I => \N__50421\
        );

    \I__12084\ : ClkMux
    port map (
            O => \N__50827\,
            I => \N__50421\
        );

    \I__12083\ : ClkMux
    port map (
            O => \N__50826\,
            I => \N__50421\
        );

    \I__12082\ : ClkMux
    port map (
            O => \N__50825\,
            I => \N__50421\
        );

    \I__12081\ : ClkMux
    port map (
            O => \N__50824\,
            I => \N__50421\
        );

    \I__12080\ : ClkMux
    port map (
            O => \N__50823\,
            I => \N__50421\
        );

    \I__12079\ : ClkMux
    port map (
            O => \N__50822\,
            I => \N__50421\
        );

    \I__12078\ : ClkMux
    port map (
            O => \N__50821\,
            I => \N__50421\
        );

    \I__12077\ : ClkMux
    port map (
            O => \N__50820\,
            I => \N__50421\
        );

    \I__12076\ : ClkMux
    port map (
            O => \N__50819\,
            I => \N__50421\
        );

    \I__12075\ : ClkMux
    port map (
            O => \N__50818\,
            I => \N__50421\
        );

    \I__12074\ : ClkMux
    port map (
            O => \N__50817\,
            I => \N__50421\
        );

    \I__12073\ : ClkMux
    port map (
            O => \N__50816\,
            I => \N__50421\
        );

    \I__12072\ : ClkMux
    port map (
            O => \N__50815\,
            I => \N__50421\
        );

    \I__12071\ : ClkMux
    port map (
            O => \N__50814\,
            I => \N__50421\
        );

    \I__12070\ : ClkMux
    port map (
            O => \N__50813\,
            I => \N__50421\
        );

    \I__12069\ : ClkMux
    port map (
            O => \N__50812\,
            I => \N__50421\
        );

    \I__12068\ : ClkMux
    port map (
            O => \N__50811\,
            I => \N__50421\
        );

    \I__12067\ : ClkMux
    port map (
            O => \N__50810\,
            I => \N__50421\
        );

    \I__12066\ : ClkMux
    port map (
            O => \N__50809\,
            I => \N__50421\
        );

    \I__12065\ : ClkMux
    port map (
            O => \N__50808\,
            I => \N__50421\
        );

    \I__12064\ : ClkMux
    port map (
            O => \N__50807\,
            I => \N__50421\
        );

    \I__12063\ : ClkMux
    port map (
            O => \N__50806\,
            I => \N__50421\
        );

    \I__12062\ : ClkMux
    port map (
            O => \N__50805\,
            I => \N__50421\
        );

    \I__12061\ : ClkMux
    port map (
            O => \N__50804\,
            I => \N__50421\
        );

    \I__12060\ : ClkMux
    port map (
            O => \N__50803\,
            I => \N__50421\
        );

    \I__12059\ : ClkMux
    port map (
            O => \N__50802\,
            I => \N__50421\
        );

    \I__12058\ : ClkMux
    port map (
            O => \N__50801\,
            I => \N__50421\
        );

    \I__12057\ : ClkMux
    port map (
            O => \N__50800\,
            I => \N__50421\
        );

    \I__12056\ : ClkMux
    port map (
            O => \N__50799\,
            I => \N__50421\
        );

    \I__12055\ : ClkMux
    port map (
            O => \N__50798\,
            I => \N__50421\
        );

    \I__12054\ : ClkMux
    port map (
            O => \N__50797\,
            I => \N__50421\
        );

    \I__12053\ : ClkMux
    port map (
            O => \N__50796\,
            I => \N__50421\
        );

    \I__12052\ : ClkMux
    port map (
            O => \N__50795\,
            I => \N__50421\
        );

    \I__12051\ : ClkMux
    port map (
            O => \N__50794\,
            I => \N__50421\
        );

    \I__12050\ : ClkMux
    port map (
            O => \N__50793\,
            I => \N__50421\
        );

    \I__12049\ : ClkMux
    port map (
            O => \N__50792\,
            I => \N__50421\
        );

    \I__12048\ : ClkMux
    port map (
            O => \N__50791\,
            I => \N__50421\
        );

    \I__12047\ : ClkMux
    port map (
            O => \N__50790\,
            I => \N__50421\
        );

    \I__12046\ : ClkMux
    port map (
            O => \N__50789\,
            I => \N__50421\
        );

    \I__12045\ : ClkMux
    port map (
            O => \N__50788\,
            I => \N__50421\
        );

    \I__12044\ : ClkMux
    port map (
            O => \N__50787\,
            I => \N__50421\
        );

    \I__12043\ : ClkMux
    port map (
            O => \N__50786\,
            I => \N__50421\
        );

    \I__12042\ : ClkMux
    port map (
            O => \N__50785\,
            I => \N__50421\
        );

    \I__12041\ : ClkMux
    port map (
            O => \N__50784\,
            I => \N__50421\
        );

    \I__12040\ : ClkMux
    port map (
            O => \N__50783\,
            I => \N__50421\
        );

    \I__12039\ : ClkMux
    port map (
            O => \N__50782\,
            I => \N__50421\
        );

    \I__12038\ : ClkMux
    port map (
            O => \N__50781\,
            I => \N__50421\
        );

    \I__12037\ : ClkMux
    port map (
            O => \N__50780\,
            I => \N__50421\
        );

    \I__12036\ : ClkMux
    port map (
            O => \N__50779\,
            I => \N__50421\
        );

    \I__12035\ : ClkMux
    port map (
            O => \N__50778\,
            I => \N__50421\
        );

    \I__12034\ : ClkMux
    port map (
            O => \N__50777\,
            I => \N__50421\
        );

    \I__12033\ : ClkMux
    port map (
            O => \N__50776\,
            I => \N__50421\
        );

    \I__12032\ : ClkMux
    port map (
            O => \N__50775\,
            I => \N__50421\
        );

    \I__12031\ : ClkMux
    port map (
            O => \N__50774\,
            I => \N__50421\
        );

    \I__12030\ : ClkMux
    port map (
            O => \N__50773\,
            I => \N__50421\
        );

    \I__12029\ : ClkMux
    port map (
            O => \N__50772\,
            I => \N__50421\
        );

    \I__12028\ : ClkMux
    port map (
            O => \N__50771\,
            I => \N__50421\
        );

    \I__12027\ : ClkMux
    port map (
            O => \N__50770\,
            I => \N__50421\
        );

    \I__12026\ : ClkMux
    port map (
            O => \N__50769\,
            I => \N__50421\
        );

    \I__12025\ : ClkMux
    port map (
            O => \N__50768\,
            I => \N__50421\
        );

    \I__12024\ : ClkMux
    port map (
            O => \N__50767\,
            I => \N__50421\
        );

    \I__12023\ : ClkMux
    port map (
            O => \N__50766\,
            I => \N__50421\
        );

    \I__12022\ : ClkMux
    port map (
            O => \N__50765\,
            I => \N__50421\
        );

    \I__12021\ : ClkMux
    port map (
            O => \N__50764\,
            I => \N__50421\
        );

    \I__12020\ : ClkMux
    port map (
            O => \N__50763\,
            I => \N__50421\
        );

    \I__12019\ : ClkMux
    port map (
            O => \N__50762\,
            I => \N__50421\
        );

    \I__12018\ : ClkMux
    port map (
            O => \N__50761\,
            I => \N__50421\
        );

    \I__12017\ : ClkMux
    port map (
            O => \N__50760\,
            I => \N__50421\
        );

    \I__12016\ : ClkMux
    port map (
            O => \N__50759\,
            I => \N__50421\
        );

    \I__12015\ : ClkMux
    port map (
            O => \N__50758\,
            I => \N__50421\
        );

    \I__12014\ : ClkMux
    port map (
            O => \N__50757\,
            I => \N__50421\
        );

    \I__12013\ : ClkMux
    port map (
            O => \N__50756\,
            I => \N__50421\
        );

    \I__12012\ : Glb2LocalMux
    port map (
            O => \N__50753\,
            I => \N__50421\
        );

    \I__12011\ : ClkMux
    port map (
            O => \N__50752\,
            I => \N__50421\
        );

    \I__12010\ : ClkMux
    port map (
            O => \N__50751\,
            I => \N__50421\
        );

    \I__12009\ : ClkMux
    port map (
            O => \N__50750\,
            I => \N__50421\
        );

    \I__12008\ : GlobalMux
    port map (
            O => \N__50421\,
            I => clock_output_0
        );

    \I__12007\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50412\
        );

    \I__12006\ : InMux
    port map (
            O => \N__50417\,
            I => \N__50407\
        );

    \I__12005\ : InMux
    port map (
            O => \N__50416\,
            I => \N__50407\
        );

    \I__12004\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50404\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__50412\,
            I => \N__50401\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50407\,
            I => \N__50398\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__50404\,
            I => \N__50395\
        );

    \I__12000\ : Glb2LocalMux
    port map (
            O => \N__50401\,
            I => \N__49890\
        );

    \I__11999\ : Glb2LocalMux
    port map (
            O => \N__50398\,
            I => \N__49890\
        );

    \I__11998\ : Glb2LocalMux
    port map (
            O => \N__50395\,
            I => \N__49890\
        );

    \I__11997\ : SRMux
    port map (
            O => \N__50394\,
            I => \N__49890\
        );

    \I__11996\ : SRMux
    port map (
            O => \N__50393\,
            I => \N__49890\
        );

    \I__11995\ : SRMux
    port map (
            O => \N__50392\,
            I => \N__49890\
        );

    \I__11994\ : SRMux
    port map (
            O => \N__50391\,
            I => \N__49890\
        );

    \I__11993\ : SRMux
    port map (
            O => \N__50390\,
            I => \N__49890\
        );

    \I__11992\ : SRMux
    port map (
            O => \N__50389\,
            I => \N__49890\
        );

    \I__11991\ : SRMux
    port map (
            O => \N__50388\,
            I => \N__49890\
        );

    \I__11990\ : SRMux
    port map (
            O => \N__50387\,
            I => \N__49890\
        );

    \I__11989\ : SRMux
    port map (
            O => \N__50386\,
            I => \N__49890\
        );

    \I__11988\ : SRMux
    port map (
            O => \N__50385\,
            I => \N__49890\
        );

    \I__11987\ : SRMux
    port map (
            O => \N__50384\,
            I => \N__49890\
        );

    \I__11986\ : SRMux
    port map (
            O => \N__50383\,
            I => \N__49890\
        );

    \I__11985\ : SRMux
    port map (
            O => \N__50382\,
            I => \N__49890\
        );

    \I__11984\ : SRMux
    port map (
            O => \N__50381\,
            I => \N__49890\
        );

    \I__11983\ : SRMux
    port map (
            O => \N__50380\,
            I => \N__49890\
        );

    \I__11982\ : SRMux
    port map (
            O => \N__50379\,
            I => \N__49890\
        );

    \I__11981\ : SRMux
    port map (
            O => \N__50378\,
            I => \N__49890\
        );

    \I__11980\ : SRMux
    port map (
            O => \N__50377\,
            I => \N__49890\
        );

    \I__11979\ : SRMux
    port map (
            O => \N__50376\,
            I => \N__49890\
        );

    \I__11978\ : SRMux
    port map (
            O => \N__50375\,
            I => \N__49890\
        );

    \I__11977\ : SRMux
    port map (
            O => \N__50374\,
            I => \N__49890\
        );

    \I__11976\ : SRMux
    port map (
            O => \N__50373\,
            I => \N__49890\
        );

    \I__11975\ : SRMux
    port map (
            O => \N__50372\,
            I => \N__49890\
        );

    \I__11974\ : SRMux
    port map (
            O => \N__50371\,
            I => \N__49890\
        );

    \I__11973\ : SRMux
    port map (
            O => \N__50370\,
            I => \N__49890\
        );

    \I__11972\ : SRMux
    port map (
            O => \N__50369\,
            I => \N__49890\
        );

    \I__11971\ : SRMux
    port map (
            O => \N__50368\,
            I => \N__49890\
        );

    \I__11970\ : SRMux
    port map (
            O => \N__50367\,
            I => \N__49890\
        );

    \I__11969\ : SRMux
    port map (
            O => \N__50366\,
            I => \N__49890\
        );

    \I__11968\ : SRMux
    port map (
            O => \N__50365\,
            I => \N__49890\
        );

    \I__11967\ : SRMux
    port map (
            O => \N__50364\,
            I => \N__49890\
        );

    \I__11966\ : SRMux
    port map (
            O => \N__50363\,
            I => \N__49890\
        );

    \I__11965\ : SRMux
    port map (
            O => \N__50362\,
            I => \N__49890\
        );

    \I__11964\ : SRMux
    port map (
            O => \N__50361\,
            I => \N__49890\
        );

    \I__11963\ : SRMux
    port map (
            O => \N__50360\,
            I => \N__49890\
        );

    \I__11962\ : SRMux
    port map (
            O => \N__50359\,
            I => \N__49890\
        );

    \I__11961\ : SRMux
    port map (
            O => \N__50358\,
            I => \N__49890\
        );

    \I__11960\ : SRMux
    port map (
            O => \N__50357\,
            I => \N__49890\
        );

    \I__11959\ : SRMux
    port map (
            O => \N__50356\,
            I => \N__49890\
        );

    \I__11958\ : SRMux
    port map (
            O => \N__50355\,
            I => \N__49890\
        );

    \I__11957\ : SRMux
    port map (
            O => \N__50354\,
            I => \N__49890\
        );

    \I__11956\ : SRMux
    port map (
            O => \N__50353\,
            I => \N__49890\
        );

    \I__11955\ : SRMux
    port map (
            O => \N__50352\,
            I => \N__49890\
        );

    \I__11954\ : SRMux
    port map (
            O => \N__50351\,
            I => \N__49890\
        );

    \I__11953\ : SRMux
    port map (
            O => \N__50350\,
            I => \N__49890\
        );

    \I__11952\ : SRMux
    port map (
            O => \N__50349\,
            I => \N__49890\
        );

    \I__11951\ : SRMux
    port map (
            O => \N__50348\,
            I => \N__49890\
        );

    \I__11950\ : SRMux
    port map (
            O => \N__50347\,
            I => \N__49890\
        );

    \I__11949\ : SRMux
    port map (
            O => \N__50346\,
            I => \N__49890\
        );

    \I__11948\ : SRMux
    port map (
            O => \N__50345\,
            I => \N__49890\
        );

    \I__11947\ : SRMux
    port map (
            O => \N__50344\,
            I => \N__49890\
        );

    \I__11946\ : SRMux
    port map (
            O => \N__50343\,
            I => \N__49890\
        );

    \I__11945\ : SRMux
    port map (
            O => \N__50342\,
            I => \N__49890\
        );

    \I__11944\ : SRMux
    port map (
            O => \N__50341\,
            I => \N__49890\
        );

    \I__11943\ : SRMux
    port map (
            O => \N__50340\,
            I => \N__49890\
        );

    \I__11942\ : SRMux
    port map (
            O => \N__50339\,
            I => \N__49890\
        );

    \I__11941\ : SRMux
    port map (
            O => \N__50338\,
            I => \N__49890\
        );

    \I__11940\ : SRMux
    port map (
            O => \N__50337\,
            I => \N__49890\
        );

    \I__11939\ : SRMux
    port map (
            O => \N__50336\,
            I => \N__49890\
        );

    \I__11938\ : SRMux
    port map (
            O => \N__50335\,
            I => \N__49890\
        );

    \I__11937\ : SRMux
    port map (
            O => \N__50334\,
            I => \N__49890\
        );

    \I__11936\ : SRMux
    port map (
            O => \N__50333\,
            I => \N__49890\
        );

    \I__11935\ : SRMux
    port map (
            O => \N__50332\,
            I => \N__49890\
        );

    \I__11934\ : SRMux
    port map (
            O => \N__50331\,
            I => \N__49890\
        );

    \I__11933\ : SRMux
    port map (
            O => \N__50330\,
            I => \N__49890\
        );

    \I__11932\ : SRMux
    port map (
            O => \N__50329\,
            I => \N__49890\
        );

    \I__11931\ : SRMux
    port map (
            O => \N__50328\,
            I => \N__49890\
        );

    \I__11930\ : SRMux
    port map (
            O => \N__50327\,
            I => \N__49890\
        );

    \I__11929\ : SRMux
    port map (
            O => \N__50326\,
            I => \N__49890\
        );

    \I__11928\ : SRMux
    port map (
            O => \N__50325\,
            I => \N__49890\
        );

    \I__11927\ : SRMux
    port map (
            O => \N__50324\,
            I => \N__49890\
        );

    \I__11926\ : SRMux
    port map (
            O => \N__50323\,
            I => \N__49890\
        );

    \I__11925\ : SRMux
    port map (
            O => \N__50322\,
            I => \N__49890\
        );

    \I__11924\ : SRMux
    port map (
            O => \N__50321\,
            I => \N__49890\
        );

    \I__11923\ : SRMux
    port map (
            O => \N__50320\,
            I => \N__49890\
        );

    \I__11922\ : SRMux
    port map (
            O => \N__50319\,
            I => \N__49890\
        );

    \I__11921\ : SRMux
    port map (
            O => \N__50318\,
            I => \N__49890\
        );

    \I__11920\ : SRMux
    port map (
            O => \N__50317\,
            I => \N__49890\
        );

    \I__11919\ : SRMux
    port map (
            O => \N__50316\,
            I => \N__49890\
        );

    \I__11918\ : SRMux
    port map (
            O => \N__50315\,
            I => \N__49890\
        );

    \I__11917\ : SRMux
    port map (
            O => \N__50314\,
            I => \N__49890\
        );

    \I__11916\ : SRMux
    port map (
            O => \N__50313\,
            I => \N__49890\
        );

    \I__11915\ : SRMux
    port map (
            O => \N__50312\,
            I => \N__49890\
        );

    \I__11914\ : SRMux
    port map (
            O => \N__50311\,
            I => \N__49890\
        );

    \I__11913\ : SRMux
    port map (
            O => \N__50310\,
            I => \N__49890\
        );

    \I__11912\ : SRMux
    port map (
            O => \N__50309\,
            I => \N__49890\
        );

    \I__11911\ : SRMux
    port map (
            O => \N__50308\,
            I => \N__49890\
        );

    \I__11910\ : SRMux
    port map (
            O => \N__50307\,
            I => \N__49890\
        );

    \I__11909\ : SRMux
    port map (
            O => \N__50306\,
            I => \N__49890\
        );

    \I__11908\ : SRMux
    port map (
            O => \N__50305\,
            I => \N__49890\
        );

    \I__11907\ : SRMux
    port map (
            O => \N__50304\,
            I => \N__49890\
        );

    \I__11906\ : SRMux
    port map (
            O => \N__50303\,
            I => \N__49890\
        );

    \I__11905\ : SRMux
    port map (
            O => \N__50302\,
            I => \N__49890\
        );

    \I__11904\ : SRMux
    port map (
            O => \N__50301\,
            I => \N__49890\
        );

    \I__11903\ : SRMux
    port map (
            O => \N__50300\,
            I => \N__49890\
        );

    \I__11902\ : SRMux
    port map (
            O => \N__50299\,
            I => \N__49890\
        );

    \I__11901\ : SRMux
    port map (
            O => \N__50298\,
            I => \N__49890\
        );

    \I__11900\ : SRMux
    port map (
            O => \N__50297\,
            I => \N__49890\
        );

    \I__11899\ : SRMux
    port map (
            O => \N__50296\,
            I => \N__49890\
        );

    \I__11898\ : SRMux
    port map (
            O => \N__50295\,
            I => \N__49890\
        );

    \I__11897\ : SRMux
    port map (
            O => \N__50294\,
            I => \N__49890\
        );

    \I__11896\ : SRMux
    port map (
            O => \N__50293\,
            I => \N__49890\
        );

    \I__11895\ : SRMux
    port map (
            O => \N__50292\,
            I => \N__49890\
        );

    \I__11894\ : SRMux
    port map (
            O => \N__50291\,
            I => \N__49890\
        );

    \I__11893\ : SRMux
    port map (
            O => \N__50290\,
            I => \N__49890\
        );

    \I__11892\ : SRMux
    port map (
            O => \N__50289\,
            I => \N__49890\
        );

    \I__11891\ : SRMux
    port map (
            O => \N__50288\,
            I => \N__49890\
        );

    \I__11890\ : SRMux
    port map (
            O => \N__50287\,
            I => \N__49890\
        );

    \I__11889\ : SRMux
    port map (
            O => \N__50286\,
            I => \N__49890\
        );

    \I__11888\ : SRMux
    port map (
            O => \N__50285\,
            I => \N__49890\
        );

    \I__11887\ : SRMux
    port map (
            O => \N__50284\,
            I => \N__49890\
        );

    \I__11886\ : SRMux
    port map (
            O => \N__50283\,
            I => \N__49890\
        );

    \I__11885\ : SRMux
    port map (
            O => \N__50282\,
            I => \N__49890\
        );

    \I__11884\ : SRMux
    port map (
            O => \N__50281\,
            I => \N__49890\
        );

    \I__11883\ : SRMux
    port map (
            O => \N__50280\,
            I => \N__49890\
        );

    \I__11882\ : SRMux
    port map (
            O => \N__50279\,
            I => \N__49890\
        );

    \I__11881\ : SRMux
    port map (
            O => \N__50278\,
            I => \N__49890\
        );

    \I__11880\ : SRMux
    port map (
            O => \N__50277\,
            I => \N__49890\
        );

    \I__11879\ : SRMux
    port map (
            O => \N__50276\,
            I => \N__49890\
        );

    \I__11878\ : SRMux
    port map (
            O => \N__50275\,
            I => \N__49890\
        );

    \I__11877\ : SRMux
    port map (
            O => \N__50274\,
            I => \N__49890\
        );

    \I__11876\ : SRMux
    port map (
            O => \N__50273\,
            I => \N__49890\
        );

    \I__11875\ : SRMux
    port map (
            O => \N__50272\,
            I => \N__49890\
        );

    \I__11874\ : SRMux
    port map (
            O => \N__50271\,
            I => \N__49890\
        );

    \I__11873\ : SRMux
    port map (
            O => \N__50270\,
            I => \N__49890\
        );

    \I__11872\ : SRMux
    port map (
            O => \N__50269\,
            I => \N__49890\
        );

    \I__11871\ : SRMux
    port map (
            O => \N__50268\,
            I => \N__49890\
        );

    \I__11870\ : SRMux
    port map (
            O => \N__50267\,
            I => \N__49890\
        );

    \I__11869\ : SRMux
    port map (
            O => \N__50266\,
            I => \N__49890\
        );

    \I__11868\ : SRMux
    port map (
            O => \N__50265\,
            I => \N__49890\
        );

    \I__11867\ : SRMux
    port map (
            O => \N__50264\,
            I => \N__49890\
        );

    \I__11866\ : SRMux
    port map (
            O => \N__50263\,
            I => \N__49890\
        );

    \I__11865\ : SRMux
    port map (
            O => \N__50262\,
            I => \N__49890\
        );

    \I__11864\ : SRMux
    port map (
            O => \N__50261\,
            I => \N__49890\
        );

    \I__11863\ : SRMux
    port map (
            O => \N__50260\,
            I => \N__49890\
        );

    \I__11862\ : SRMux
    port map (
            O => \N__50259\,
            I => \N__49890\
        );

    \I__11861\ : SRMux
    port map (
            O => \N__50258\,
            I => \N__49890\
        );

    \I__11860\ : SRMux
    port map (
            O => \N__50257\,
            I => \N__49890\
        );

    \I__11859\ : SRMux
    port map (
            O => \N__50256\,
            I => \N__49890\
        );

    \I__11858\ : SRMux
    port map (
            O => \N__50255\,
            I => \N__49890\
        );

    \I__11857\ : SRMux
    port map (
            O => \N__50254\,
            I => \N__49890\
        );

    \I__11856\ : SRMux
    port map (
            O => \N__50253\,
            I => \N__49890\
        );

    \I__11855\ : SRMux
    port map (
            O => \N__50252\,
            I => \N__49890\
        );

    \I__11854\ : SRMux
    port map (
            O => \N__50251\,
            I => \N__49890\
        );

    \I__11853\ : SRMux
    port map (
            O => \N__50250\,
            I => \N__49890\
        );

    \I__11852\ : SRMux
    port map (
            O => \N__50249\,
            I => \N__49890\
        );

    \I__11851\ : SRMux
    port map (
            O => \N__50248\,
            I => \N__49890\
        );

    \I__11850\ : SRMux
    port map (
            O => \N__50247\,
            I => \N__49890\
        );

    \I__11849\ : SRMux
    port map (
            O => \N__50246\,
            I => \N__49890\
        );

    \I__11848\ : SRMux
    port map (
            O => \N__50245\,
            I => \N__49890\
        );

    \I__11847\ : SRMux
    port map (
            O => \N__50244\,
            I => \N__49890\
        );

    \I__11846\ : SRMux
    port map (
            O => \N__50243\,
            I => \N__49890\
        );

    \I__11845\ : SRMux
    port map (
            O => \N__50242\,
            I => \N__49890\
        );

    \I__11844\ : SRMux
    port map (
            O => \N__50241\,
            I => \N__49890\
        );

    \I__11843\ : SRMux
    port map (
            O => \N__50240\,
            I => \N__49890\
        );

    \I__11842\ : SRMux
    port map (
            O => \N__50239\,
            I => \N__49890\
        );

    \I__11841\ : SRMux
    port map (
            O => \N__50238\,
            I => \N__49890\
        );

    \I__11840\ : SRMux
    port map (
            O => \N__50237\,
            I => \N__49890\
        );

    \I__11839\ : SRMux
    port map (
            O => \N__50236\,
            I => \N__49890\
        );

    \I__11838\ : SRMux
    port map (
            O => \N__50235\,
            I => \N__49890\
        );

    \I__11837\ : SRMux
    port map (
            O => \N__50234\,
            I => \N__49890\
        );

    \I__11836\ : SRMux
    port map (
            O => \N__50233\,
            I => \N__49890\
        );

    \I__11835\ : SRMux
    port map (
            O => \N__50232\,
            I => \N__49890\
        );

    \I__11834\ : SRMux
    port map (
            O => \N__50231\,
            I => \N__49890\
        );

    \I__11833\ : SRMux
    port map (
            O => \N__50230\,
            I => \N__49890\
        );

    \I__11832\ : SRMux
    port map (
            O => \N__50229\,
            I => \N__49890\
        );

    \I__11831\ : GlobalMux
    port map (
            O => \N__49890\,
            I => \N__49887\
        );

    \I__11830\ : gio2CtrlBuf
    port map (
            O => \N__49887\,
            I => red_c_g
        );

    \I__11829\ : InMux
    port map (
            O => \N__49884\,
            I => \N__49879\
        );

    \I__11828\ : InMux
    port map (
            O => \N__49883\,
            I => \N__49876\
        );

    \I__11827\ : InMux
    port map (
            O => \N__49882\,
            I => \N__49873\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__49879\,
            I => \N__49858\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__49876\,
            I => \N__49858\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__49873\,
            I => \N__49858\
        );

    \I__11823\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49855\
        );

    \I__11822\ : InMux
    port map (
            O => \N__49871\,
            I => \N__49848\
        );

    \I__11821\ : InMux
    port map (
            O => \N__49870\,
            I => \N__49848\
        );

    \I__11820\ : InMux
    port map (
            O => \N__49869\,
            I => \N__49848\
        );

    \I__11819\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49839\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49839\
        );

    \I__11817\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49839\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49865\,
            I => \N__49839\
        );

    \I__11815\ : Span4Mux_s3_v
    port map (
            O => \N__49858\,
            I => \N__49830\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__49855\,
            I => \N__49830\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__49848\,
            I => \N__49830\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__49839\,
            I => \N__49830\
        );

    \I__11811\ : Span4Mux_v
    port map (
            O => \N__49830\,
            I => \N__49827\
        );

    \I__11810\ : Span4Mux_v
    port map (
            O => \N__49827\,
            I => \N__49822\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49826\,
            I => \N__49819\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49811\
        );

    \I__11807\ : Span4Mux_v
    port map (
            O => \N__49822\,
            I => \N__49806\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__49819\,
            I => \N__49806\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49801\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49817\,
            I => \N__49801\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49816\,
            I => \N__49798\
        );

    \I__11802\ : CascadeMux
    port map (
            O => \N__49815\,
            I => \N__49786\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49814\,
            I => \N__49766\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__49811\,
            I => \N__49763\
        );

    \I__11799\ : Span4Mux_v
    port map (
            O => \N__49806\,
            I => \N__49756\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__49801\,
            I => \N__49756\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__49798\,
            I => \N__49756\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49797\,
            I => \N__49753\
        );

    \I__11795\ : InMux
    port map (
            O => \N__49796\,
            I => \N__49746\
        );

    \I__11794\ : InMux
    port map (
            O => \N__49795\,
            I => \N__49746\
        );

    \I__11793\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49746\
        );

    \I__11792\ : InMux
    port map (
            O => \N__49793\,
            I => \N__49737\
        );

    \I__11791\ : InMux
    port map (
            O => \N__49792\,
            I => \N__49737\
        );

    \I__11790\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49737\
        );

    \I__11789\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49737\
        );

    \I__11788\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49730\
        );

    \I__11787\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49730\
        );

    \I__11786\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49730\
        );

    \I__11785\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49727\
        );

    \I__11784\ : CascadeMux
    port map (
            O => \N__49783\,
            I => \N__49723\
        );

    \I__11783\ : CascadeMux
    port map (
            O => \N__49782\,
            I => \N__49719\
        );

    \I__11782\ : CascadeMux
    port map (
            O => \N__49781\,
            I => \N__49715\
        );

    \I__11781\ : CascadeMux
    port map (
            O => \N__49780\,
            I => \N__49711\
        );

    \I__11780\ : CascadeMux
    port map (
            O => \N__49779\,
            I => \N__49707\
        );

    \I__11779\ : CascadeMux
    port map (
            O => \N__49778\,
            I => \N__49703\
        );

    \I__11778\ : CascadeMux
    port map (
            O => \N__49777\,
            I => \N__49699\
        );

    \I__11777\ : CascadeMux
    port map (
            O => \N__49776\,
            I => \N__49695\
        );

    \I__11776\ : CascadeMux
    port map (
            O => \N__49775\,
            I => \N__49692\
        );

    \I__11775\ : CascadeMux
    port map (
            O => \N__49774\,
            I => \N__49688\
        );

    \I__11774\ : CascadeMux
    port map (
            O => \N__49773\,
            I => \N__49684\
        );

    \I__11773\ : CascadeMux
    port map (
            O => \N__49772\,
            I => \N__49680\
        );

    \I__11772\ : CascadeMux
    port map (
            O => \N__49771\,
            I => \N__49675\
        );

    \I__11771\ : CascadeMux
    port map (
            O => \N__49770\,
            I => \N__49671\
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__49769\,
            I => \N__49667\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__49766\,
            I => \N__49661\
        );

    \I__11768\ : Span4Mux_v
    port map (
            O => \N__49763\,
            I => \N__49661\
        );

    \I__11767\ : Span4Mux_v
    port map (
            O => \N__49756\,
            I => \N__49649\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__49753\,
            I => \N__49649\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__49746\,
            I => \N__49649\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49737\,
            I => \N__49649\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__49730\,
            I => \N__49646\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__49727\,
            I => \N__49643\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49726\,
            I => \N__49640\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49625\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49722\,
            I => \N__49625\
        );

    \I__11758\ : InMux
    port map (
            O => \N__49719\,
            I => \N__49625\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49718\,
            I => \N__49625\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49715\,
            I => \N__49625\
        );

    \I__11755\ : InMux
    port map (
            O => \N__49714\,
            I => \N__49625\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49711\,
            I => \N__49625\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49608\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49707\,
            I => \N__49608\
        );

    \I__11751\ : InMux
    port map (
            O => \N__49706\,
            I => \N__49608\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49703\,
            I => \N__49608\
        );

    \I__11749\ : InMux
    port map (
            O => \N__49702\,
            I => \N__49608\
        );

    \I__11748\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49608\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49608\
        );

    \I__11746\ : InMux
    port map (
            O => \N__49695\,
            I => \N__49608\
        );

    \I__11745\ : InMux
    port map (
            O => \N__49692\,
            I => \N__49591\
        );

    \I__11744\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49591\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49688\,
            I => \N__49591\
        );

    \I__11742\ : InMux
    port map (
            O => \N__49687\,
            I => \N__49591\
        );

    \I__11741\ : InMux
    port map (
            O => \N__49684\,
            I => \N__49591\
        );

    \I__11740\ : InMux
    port map (
            O => \N__49683\,
            I => \N__49591\
        );

    \I__11739\ : InMux
    port map (
            O => \N__49680\,
            I => \N__49591\
        );

    \I__11738\ : InMux
    port map (
            O => \N__49679\,
            I => \N__49591\
        );

    \I__11737\ : InMux
    port map (
            O => \N__49678\,
            I => \N__49576\
        );

    \I__11736\ : InMux
    port map (
            O => \N__49675\,
            I => \N__49576\
        );

    \I__11735\ : InMux
    port map (
            O => \N__49674\,
            I => \N__49576\
        );

    \I__11734\ : InMux
    port map (
            O => \N__49671\,
            I => \N__49576\
        );

    \I__11733\ : InMux
    port map (
            O => \N__49670\,
            I => \N__49576\
        );

    \I__11732\ : InMux
    port map (
            O => \N__49667\,
            I => \N__49576\
        );

    \I__11731\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49576\
        );

    \I__11730\ : IoSpan4Mux
    port map (
            O => \N__49661\,
            I => \N__49573\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49660\,
            I => \N__49568\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49659\,
            I => \N__49568\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49658\,
            I => \N__49565\
        );

    \I__11726\ : Span4Mux_v
    port map (
            O => \N__49649\,
            I => \N__49562\
        );

    \I__11725\ : Span4Mux_v
    port map (
            O => \N__49646\,
            I => \N__49559\
        );

    \I__11724\ : Span4Mux_v
    port map (
            O => \N__49643\,
            I => \N__49554\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__49640\,
            I => \N__49554\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49625\,
            I => \N__49545\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__49608\,
            I => \N__49545\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__49591\,
            I => \N__49545\
        );

    \I__11719\ : LocalMux
    port map (
            O => \N__49576\,
            I => \N__49545\
        );

    \I__11718\ : Span4Mux_s0_v
    port map (
            O => \N__49573\,
            I => \N__49542\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__49568\,
            I => \N__49537\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__49565\,
            I => \N__49537\
        );

    \I__11715\ : Sp12to4
    port map (
            O => \N__49562\,
            I => \N__49534\
        );

    \I__11714\ : Sp12to4
    port map (
            O => \N__49559\,
            I => \N__49531\
        );

    \I__11713\ : Span4Mux_h
    port map (
            O => \N__49554\,
            I => \N__49526\
        );

    \I__11712\ : Span4Mux_v
    port map (
            O => \N__49545\,
            I => \N__49526\
        );

    \I__11711\ : Span4Mux_v
    port map (
            O => \N__49542\,
            I => \N__49523\
        );

    \I__11710\ : Span4Mux_s3_h
    port map (
            O => \N__49537\,
            I => \N__49520\
        );

    \I__11709\ : Span12Mux_s10_h
    port map (
            O => \N__49534\,
            I => \N__49517\
        );

    \I__11708\ : Span12Mux_s10_h
    port map (
            O => \N__49531\,
            I => \N__49512\
        );

    \I__11707\ : Sp12to4
    port map (
            O => \N__49526\,
            I => \N__49512\
        );

    \I__11706\ : Sp12to4
    port map (
            O => \N__49523\,
            I => \N__49507\
        );

    \I__11705\ : Sp12to4
    port map (
            O => \N__49520\,
            I => \N__49507\
        );

    \I__11704\ : Span12Mux_h
    port map (
            O => \N__49517\,
            I => \N__49500\
        );

    \I__11703\ : Span12Mux_h
    port map (
            O => \N__49512\,
            I => \N__49500\
        );

    \I__11702\ : Span12Mux_v
    port map (
            O => \N__49507\,
            I => \N__49500\
        );

    \I__11701\ : Odrv12
    port map (
            O => \N__49500\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11700\ : InMux
    port map (
            O => \N__49497\,
            I => \N__49493\
        );

    \I__11699\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49489\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__49493\,
            I => \N__49486\
        );

    \I__11697\ : InMux
    port map (
            O => \N__49492\,
            I => \N__49483\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__49489\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__11695\ : Odrv4
    port map (
            O => \N__49486\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49483\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49476\,
            I => \N__49470\
        );

    \I__11692\ : InMux
    port map (
            O => \N__49475\,
            I => \N__49467\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49474\,
            I => \N__49464\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49473\,
            I => \N__49461\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__49470\,
            I => \N__49458\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__49467\,
            I => \N__49453\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__49464\,
            I => \N__49453\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__49461\,
            I => \N__49450\
        );

    \I__11685\ : Span4Mux_v
    port map (
            O => \N__49458\,
            I => \N__49443\
        );

    \I__11684\ : Span4Mux_v
    port map (
            O => \N__49453\,
            I => \N__49443\
        );

    \I__11683\ : Span4Mux_v
    port map (
            O => \N__49450\,
            I => \N__49443\
        );

    \I__11682\ : Odrv4
    port map (
            O => \N__49443\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__11681\ : CascadeMux
    port map (
            O => \N__49440\,
            I => \N__49436\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49439\,
            I => \N__49431\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49431\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__49431\,
            I => \N__49428\
        );

    \I__11677\ : Odrv4
    port map (
            O => \N__49428\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__11676\ : CascadeMux
    port map (
            O => \N__49425\,
            I => \N__49422\
        );

    \I__11675\ : InMux
    port map (
            O => \N__49422\,
            I => \N__49416\
        );

    \I__11674\ : InMux
    port map (
            O => \N__49421\,
            I => \N__49413\
        );

    \I__11673\ : InMux
    port map (
            O => \N__49420\,
            I => \N__49410\
        );

    \I__11672\ : InMux
    port map (
            O => \N__49419\,
            I => \N__49407\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__49416\,
            I => \N__49404\
        );

    \I__11670\ : LocalMux
    port map (
            O => \N__49413\,
            I => \N__49401\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__49410\,
            I => \N__49396\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__49407\,
            I => \N__49396\
        );

    \I__11667\ : Span4Mux_h
    port map (
            O => \N__49404\,
            I => \N__49393\
        );

    \I__11666\ : Span4Mux_v
    port map (
            O => \N__49401\,
            I => \N__49390\
        );

    \I__11665\ : Span4Mux_v
    port map (
            O => \N__49396\,
            I => \N__49385\
        );

    \I__11664\ : Span4Mux_v
    port map (
            O => \N__49393\,
            I => \N__49385\
        );

    \I__11663\ : Odrv4
    port map (
            O => \N__49390\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__49385\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49380\,
            I => \N__49377\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__49377\,
            I => \N__49374\
        );

    \I__11659\ : Span4Mux_h
    port map (
            O => \N__49374\,
            I => \N__49369\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49373\,
            I => \N__49366\
        );

    \I__11657\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49363\
        );

    \I__11656\ : Span4Mux_v
    port map (
            O => \N__49369\,
            I => \N__49360\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__49366\,
            I => \N__49357\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__49363\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__11653\ : Odrv4
    port map (
            O => \N__49360\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__11652\ : Odrv4
    port map (
            O => \N__49357\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49347\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__49347\,
            I => \N__49344\
        );

    \I__11649\ : Odrv4
    port map (
            O => \N__49344\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__11648\ : CascadeMux
    port map (
            O => \N__49341\,
            I => \N__49338\
        );

    \I__11647\ : InMux
    port map (
            O => \N__49338\,
            I => \N__49332\
        );

    \I__11646\ : InMux
    port map (
            O => \N__49337\,
            I => \N__49332\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__49332\,
            I => \N__49329\
        );

    \I__11644\ : Span4Mux_h
    port map (
            O => \N__49329\,
            I => \N__49326\
        );

    \I__11643\ : Odrv4
    port map (
            O => \N__49326\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__11642\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49319\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49315\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__49319\,
            I => \N__49312\
        );

    \I__11639\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49309\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__49315\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__11637\ : Odrv12
    port map (
            O => \N__49312\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__11636\ : LocalMux
    port map (
            O => \N__49309\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49298\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49293\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__49298\,
            I => \N__49290\
        );

    \I__11632\ : InMux
    port map (
            O => \N__49297\,
            I => \N__49285\
        );

    \I__11631\ : InMux
    port map (
            O => \N__49296\,
            I => \N__49285\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__49293\,
            I => \N__49282\
        );

    \I__11629\ : Span4Mux_h
    port map (
            O => \N__49290\,
            I => \N__49279\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__49285\,
            I => \N__49276\
        );

    \I__11627\ : Span4Mux_h
    port map (
            O => \N__49282\,
            I => \N__49271\
        );

    \I__11626\ : Span4Mux_v
    port map (
            O => \N__49279\,
            I => \N__49271\
        );

    \I__11625\ : Span4Mux_h
    port map (
            O => \N__49276\,
            I => \N__49268\
        );

    \I__11624\ : Odrv4
    port map (
            O => \N__49271\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__11623\ : Odrv4
    port map (
            O => \N__49268\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__11622\ : InMux
    port map (
            O => \N__49263\,
            I => \N__49260\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__49260\,
            I => \N__49257\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__49257\,
            I => \N__49254\
        );

    \I__11619\ : Odrv4
    port map (
            O => \N__49254\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__11618\ : CEMux
    port map (
            O => \N__49251\,
            I => \N__49212\
        );

    \I__11617\ : CEMux
    port map (
            O => \N__49250\,
            I => \N__49212\
        );

    \I__11616\ : CEMux
    port map (
            O => \N__49249\,
            I => \N__49212\
        );

    \I__11615\ : CEMux
    port map (
            O => \N__49248\,
            I => \N__49212\
        );

    \I__11614\ : CEMux
    port map (
            O => \N__49247\,
            I => \N__49212\
        );

    \I__11613\ : CEMux
    port map (
            O => \N__49246\,
            I => \N__49212\
        );

    \I__11612\ : CEMux
    port map (
            O => \N__49245\,
            I => \N__49212\
        );

    \I__11611\ : CEMux
    port map (
            O => \N__49244\,
            I => \N__49212\
        );

    \I__11610\ : CEMux
    port map (
            O => \N__49243\,
            I => \N__49212\
        );

    \I__11609\ : CEMux
    port map (
            O => \N__49242\,
            I => \N__49212\
        );

    \I__11608\ : CEMux
    port map (
            O => \N__49241\,
            I => \N__49212\
        );

    \I__11607\ : CEMux
    port map (
            O => \N__49240\,
            I => \N__49212\
        );

    \I__11606\ : CEMux
    port map (
            O => \N__49239\,
            I => \N__49212\
        );

    \I__11605\ : GlobalMux
    port map (
            O => \N__49212\,
            I => \N__49209\
        );

    \I__11604\ : gio2CtrlBuf
    port map (
            O => \N__49209\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__11603\ : InMux
    port map (
            O => \N__49206\,
            I => \N__49202\
        );

    \I__11602\ : InMux
    port map (
            O => \N__49205\,
            I => \N__49197\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__49202\,
            I => \N__49194\
        );

    \I__11600\ : InMux
    port map (
            O => \N__49201\,
            I => \N__49189\
        );

    \I__11599\ : InMux
    port map (
            O => \N__49200\,
            I => \N__49189\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__49197\,
            I => \N__49186\
        );

    \I__11597\ : Span4Mux_v
    port map (
            O => \N__49194\,
            I => \N__49183\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__49189\,
            I => \N__49180\
        );

    \I__11595\ : Span4Mux_v
    port map (
            O => \N__49186\,
            I => \N__49177\
        );

    \I__11594\ : Span4Mux_v
    port map (
            O => \N__49183\,
            I => \N__49174\
        );

    \I__11593\ : Span4Mux_h
    port map (
            O => \N__49180\,
            I => \N__49171\
        );

    \I__11592\ : Odrv4
    port map (
            O => \N__49177\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__49174\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__49171\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__11589\ : InMux
    port map (
            O => \N__49164\,
            I => \N__49161\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__49161\,
            I => \N__49158\
        );

    \I__11587\ : Span4Mux_v
    port map (
            O => \N__49158\,
            I => \N__49155\
        );

    \I__11586\ : Span4Mux_v
    port map (
            O => \N__49155\,
            I => \N__49150\
        );

    \I__11585\ : InMux
    port map (
            O => \N__49154\,
            I => \N__49147\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49153\,
            I => \N__49144\
        );

    \I__11583\ : Span4Mux_h
    port map (
            O => \N__49150\,
            I => \N__49141\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__49147\,
            I => \N__49138\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__49144\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__11580\ : Odrv4
    port map (
            O => \N__49141\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__11579\ : Odrv4
    port map (
            O => \N__49138\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__11578\ : InMux
    port map (
            O => \N__49131\,
            I => \N__49127\
        );

    \I__11577\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49124\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__49127\,
            I => \N__49121\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__49124\,
            I => \N__49116\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__49121\,
            I => \N__49113\
        );

    \I__11573\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49110\
        );

    \I__11572\ : InMux
    port map (
            O => \N__49119\,
            I => \N__49107\
        );

    \I__11571\ : Span4Mux_v
    port map (
            O => \N__49116\,
            I => \N__49100\
        );

    \I__11570\ : Span4Mux_h
    port map (
            O => \N__49113\,
            I => \N__49100\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__49110\,
            I => \N__49100\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__49107\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__11567\ : Odrv4
    port map (
            O => \N__49100\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__11566\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49069\
        );

    \I__11565\ : InMux
    port map (
            O => \N__49094\,
            I => \N__49069\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49093\,
            I => \N__49060\
        );

    \I__11563\ : InMux
    port map (
            O => \N__49092\,
            I => \N__49060\
        );

    \I__11562\ : InMux
    port map (
            O => \N__49091\,
            I => \N__49060\
        );

    \I__11561\ : InMux
    port map (
            O => \N__49090\,
            I => \N__49060\
        );

    \I__11560\ : InMux
    port map (
            O => \N__49089\,
            I => \N__49051\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49088\,
            I => \N__49051\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49051\
        );

    \I__11557\ : InMux
    port map (
            O => \N__49086\,
            I => \N__49051\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49085\,
            I => \N__49042\
        );

    \I__11555\ : InMux
    port map (
            O => \N__49084\,
            I => \N__49042\
        );

    \I__11554\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49042\
        );

    \I__11553\ : InMux
    port map (
            O => \N__49082\,
            I => \N__49042\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49033\
        );

    \I__11551\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49033\
        );

    \I__11550\ : InMux
    port map (
            O => \N__49079\,
            I => \N__49033\
        );

    \I__11549\ : InMux
    port map (
            O => \N__49078\,
            I => \N__49033\
        );

    \I__11548\ : InMux
    port map (
            O => \N__49077\,
            I => \N__49016\
        );

    \I__11547\ : InMux
    port map (
            O => \N__49076\,
            I => \N__49016\
        );

    \I__11546\ : InMux
    port map (
            O => \N__49075\,
            I => \N__49016\
        );

    \I__11545\ : InMux
    port map (
            O => \N__49074\,
            I => \N__49016\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__49069\,
            I => \N__49005\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__49005\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__49051\,
            I => \N__49005\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__49042\,
            I => \N__49005\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__49033\,
            I => \N__49005\
        );

    \I__11539\ : InMux
    port map (
            O => \N__49032\,
            I => \N__48996\
        );

    \I__11538\ : InMux
    port map (
            O => \N__49031\,
            I => \N__48996\
        );

    \I__11537\ : InMux
    port map (
            O => \N__49030\,
            I => \N__48996\
        );

    \I__11536\ : InMux
    port map (
            O => \N__49029\,
            I => \N__48996\
        );

    \I__11535\ : InMux
    port map (
            O => \N__49028\,
            I => \N__48987\
        );

    \I__11534\ : InMux
    port map (
            O => \N__49027\,
            I => \N__48987\
        );

    \I__11533\ : InMux
    port map (
            O => \N__49026\,
            I => \N__48987\
        );

    \I__11532\ : InMux
    port map (
            O => \N__49025\,
            I => \N__48987\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__49016\,
            I => \N__48980\
        );

    \I__11530\ : Span4Mux_v
    port map (
            O => \N__49005\,
            I => \N__48980\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__48996\,
            I => \N__48980\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__48987\,
            I => \N__48977\
        );

    \I__11527\ : Span4Mux_h
    port map (
            O => \N__48980\,
            I => \N__48974\
        );

    \I__11526\ : Span4Mux_h
    port map (
            O => \N__48977\,
            I => \N__48971\
        );

    \I__11525\ : Span4Mux_v
    port map (
            O => \N__48974\,
            I => \N__48968\
        );

    \I__11524\ : Odrv4
    port map (
            O => \N__48971\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__11523\ : Odrv4
    port map (
            O => \N__48968\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__11522\ : InMux
    port map (
            O => \N__48963\,
            I => \N__48958\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48955\
        );

    \I__11520\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48952\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__48958\,
            I => \N__48949\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__48955\,
            I => \N__48946\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__48952\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11516\ : Odrv12
    port map (
            O => \N__48949\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11515\ : Odrv4
    port map (
            O => \N__48946\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__48939\,
            I => \N__48933\
        );

    \I__11513\ : InMux
    port map (
            O => \N__48938\,
            I => \N__48930\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48937\,
            I => \N__48927\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48924\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48921\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__48930\,
            I => \N__48918\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__48927\,
            I => \N__48915\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__48924\,
            I => \N__48912\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__48921\,
            I => \N__48909\
        );

    \I__11505\ : Span4Mux_v
    port map (
            O => \N__48918\,
            I => \N__48902\
        );

    \I__11504\ : Span4Mux_v
    port map (
            O => \N__48915\,
            I => \N__48902\
        );

    \I__11503\ : Span4Mux_v
    port map (
            O => \N__48912\,
            I => \N__48902\
        );

    \I__11502\ : Span4Mux_h
    port map (
            O => \N__48909\,
            I => \N__48899\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__48902\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__48899\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__11499\ : CascadeMux
    port map (
            O => \N__48894\,
            I => \N__48890\
        );

    \I__11498\ : CascadeMux
    port map (
            O => \N__48893\,
            I => \N__48887\
        );

    \I__11497\ : InMux
    port map (
            O => \N__48890\,
            I => \N__48882\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48882\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__48882\,
            I => \N__48879\
        );

    \I__11494\ : Odrv12
    port map (
            O => \N__48879\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__11493\ : CEMux
    port map (
            O => \N__48876\,
            I => \N__48872\
        );

    \I__11492\ : CEMux
    port map (
            O => \N__48875\,
            I => \N__48869\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__48872\,
            I => \N__48863\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__48869\,
            I => \N__48857\
        );

    \I__11489\ : CEMux
    port map (
            O => \N__48868\,
            I => \N__48854\
        );

    \I__11488\ : CEMux
    port map (
            O => \N__48867\,
            I => \N__48848\
        );

    \I__11487\ : CEMux
    port map (
            O => \N__48866\,
            I => \N__48845\
        );

    \I__11486\ : Span4Mux_h
    port map (
            O => \N__48863\,
            I => \N__48830\
        );

    \I__11485\ : CEMux
    port map (
            O => \N__48862\,
            I => \N__48827\
        );

    \I__11484\ : CEMux
    port map (
            O => \N__48861\,
            I => \N__48821\
        );

    \I__11483\ : CEMux
    port map (
            O => \N__48860\,
            I => \N__48818\
        );

    \I__11482\ : Span4Mux_v
    port map (
            O => \N__48857\,
            I => \N__48813\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__48854\,
            I => \N__48813\
        );

    \I__11480\ : CEMux
    port map (
            O => \N__48853\,
            I => \N__48806\
        );

    \I__11479\ : CEMux
    port map (
            O => \N__48852\,
            I => \N__48803\
        );

    \I__11478\ : CEMux
    port map (
            O => \N__48851\,
            I => \N__48800\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48848\,
            I => \N__48797\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__48845\,
            I => \N__48794\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48844\,
            I => \N__48787\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48843\,
            I => \N__48787\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48842\,
            I => \N__48787\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48841\,
            I => \N__48778\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48778\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48778\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48778\
        );

    \I__11468\ : CEMux
    port map (
            O => \N__48837\,
            I => \N__48775\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48836\,
            I => \N__48766\
        );

    \I__11466\ : InMux
    port map (
            O => \N__48835\,
            I => \N__48766\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48766\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48766\
        );

    \I__11463\ : Span4Mux_h
    port map (
            O => \N__48830\,
            I => \N__48761\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__48827\,
            I => \N__48761\
        );

    \I__11461\ : CEMux
    port map (
            O => \N__48826\,
            I => \N__48758\
        );

    \I__11460\ : CEMux
    port map (
            O => \N__48825\,
            I => \N__48755\
        );

    \I__11459\ : CEMux
    port map (
            O => \N__48824\,
            I => \N__48748\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__48821\,
            I => \N__48745\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__48818\,
            I => \N__48742\
        );

    \I__11456\ : Span4Mux_v
    port map (
            O => \N__48813\,
            I => \N__48739\
        );

    \I__11455\ : CEMux
    port map (
            O => \N__48812\,
            I => \N__48736\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48811\,
            I => \N__48729\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48810\,
            I => \N__48729\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48809\,
            I => \N__48729\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__48806\,
            I => \N__48724\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__48803\,
            I => \N__48724\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__48800\,
            I => \N__48708\
        );

    \I__11448\ : Span4Mux_h
    port map (
            O => \N__48797\,
            I => \N__48693\
        );

    \I__11447\ : Span4Mux_h
    port map (
            O => \N__48794\,
            I => \N__48693\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__48787\,
            I => \N__48693\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__48778\,
            I => \N__48693\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__48775\,
            I => \N__48693\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48766\,
            I => \N__48693\
        );

    \I__11442\ : Span4Mux_h
    port map (
            O => \N__48761\,
            I => \N__48693\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__48758\,
            I => \N__48690\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48755\,
            I => \N__48687\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48678\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48678\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48752\,
            I => \N__48678\
        );

    \I__11436\ : InMux
    port map (
            O => \N__48751\,
            I => \N__48678\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48748\,
            I => \N__48669\
        );

    \I__11434\ : Span4Mux_v
    port map (
            O => \N__48745\,
            I => \N__48669\
        );

    \I__11433\ : Span4Mux_h
    port map (
            O => \N__48742\,
            I => \N__48669\
        );

    \I__11432\ : Span4Mux_h
    port map (
            O => \N__48739\,
            I => \N__48669\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__48736\,
            I => \N__48666\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__48729\,
            I => \N__48661\
        );

    \I__11429\ : Span4Mux_v
    port map (
            O => \N__48724\,
            I => \N__48661\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48723\,
            I => \N__48652\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48722\,
            I => \N__48652\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48652\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48652\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48719\,
            I => \N__48643\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48643\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48643\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48716\,
            I => \N__48643\
        );

    \I__11420\ : InMux
    port map (
            O => \N__48715\,
            I => \N__48634\
        );

    \I__11419\ : InMux
    port map (
            O => \N__48714\,
            I => \N__48634\
        );

    \I__11418\ : InMux
    port map (
            O => \N__48713\,
            I => \N__48634\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48712\,
            I => \N__48634\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48711\,
            I => \N__48631\
        );

    \I__11415\ : Sp12to4
    port map (
            O => \N__48708\,
            I => \N__48628\
        );

    \I__11414\ : Span4Mux_v
    port map (
            O => \N__48693\,
            I => \N__48625\
        );

    \I__11413\ : Span4Mux_h
    port map (
            O => \N__48690\,
            I => \N__48616\
        );

    \I__11412\ : Span4Mux_v
    port map (
            O => \N__48687\,
            I => \N__48616\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48616\
        );

    \I__11410\ : Span4Mux_h
    port map (
            O => \N__48669\,
            I => \N__48616\
        );

    \I__11409\ : Odrv4
    port map (
            O => \N__48666\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11408\ : Odrv4
    port map (
            O => \N__48661\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48652\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48643\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48634\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48631\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11403\ : Odrv12
    port map (
            O => \N__48628\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__48625\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11401\ : Odrv4
    port map (
            O => \N__48616\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48597\,
            I => \N__48594\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48594\,
            I => \N__48589\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48586\
        );

    \I__11397\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48583\
        );

    \I__11396\ : Span4Mux_h
    port map (
            O => \N__48589\,
            I => \N__48578\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48586\,
            I => \N__48578\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__48583\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__11393\ : Odrv4
    port map (
            O => \N__48578\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48573\,
            I => \N__48568\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48562\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48562\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48559\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48556\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__48562\,
            I => \N__48553\
        );

    \I__11386\ : Span4Mux_h
    port map (
            O => \N__48559\,
            I => \N__48550\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__48556\,
            I => \N__48547\
        );

    \I__11384\ : Span4Mux_h
    port map (
            O => \N__48553\,
            I => \N__48544\
        );

    \I__11383\ : Odrv4
    port map (
            O => \N__48550\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__48547\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__48544\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48534\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48534\,
            I => \N__48531\
        );

    \I__11378\ : Span4Mux_v
    port map (
            O => \N__48531\,
            I => \N__48528\
        );

    \I__11377\ : Odrv4
    port map (
            O => \N__48528\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48525\,
            I => \N__48520\
        );

    \I__11375\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48517\
        );

    \I__11374\ : InMux
    port map (
            O => \N__48523\,
            I => \N__48514\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48520\,
            I => \N__48511\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48508\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__48514\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__11370\ : Odrv12
    port map (
            O => \N__48511\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__48508\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__11368\ : InMux
    port map (
            O => \N__48501\,
            I => \N__48497\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48494\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48489\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__48494\,
            I => \N__48486\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48483\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48492\,
            I => \N__48480\
        );

    \I__11362\ : Odrv12
    port map (
            O => \N__48489\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11361\ : Odrv4
    port map (
            O => \N__48486\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__48483\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__48480\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__11358\ : InMux
    port map (
            O => \N__48471\,
            I => \N__48468\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__48468\,
            I => \N__48465\
        );

    \I__11356\ : Span4Mux_v
    port map (
            O => \N__48465\,
            I => \N__48462\
        );

    \I__11355\ : Odrv4
    port map (
            O => \N__48462\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__11354\ : InMux
    port map (
            O => \N__48459\,
            I => \N__48456\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48456\,
            I => \N__48451\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48455\,
            I => \N__48448\
        );

    \I__11351\ : InMux
    port map (
            O => \N__48454\,
            I => \N__48445\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__48451\,
            I => \N__48442\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__48448\,
            I => \N__48439\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__48445\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__48442\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__11346\ : Odrv12
    port map (
            O => \N__48439\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48426\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48421\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48421\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48418\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48415\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__48421\,
            I => \N__48412\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__48418\,
            I => \N__48409\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__48415\,
            I => \N__48404\
        );

    \I__11337\ : Span4Mux_v
    port map (
            O => \N__48412\,
            I => \N__48404\
        );

    \I__11336\ : Odrv12
    port map (
            O => \N__48409\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__11335\ : Odrv4
    port map (
            O => \N__48404\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__11334\ : CascadeMux
    port map (
            O => \N__48399\,
            I => \N__48396\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48393\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__48393\,
            I => \N__48390\
        );

    \I__11331\ : Span4Mux_v
    port map (
            O => \N__48390\,
            I => \N__48387\
        );

    \I__11330\ : Odrv4
    port map (
            O => \N__48387\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__11329\ : CascadeMux
    port map (
            O => \N__48384\,
            I => \N__48378\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48373\
        );

    \I__11327\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48373\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48381\,
            I => \N__48370\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48378\,
            I => \N__48367\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48364\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__48370\,
            I => \N__48361\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48358\
        );

    \I__11321\ : Span4Mux_h
    port map (
            O => \N__48364\,
            I => \N__48355\
        );

    \I__11320\ : Span4Mux_h
    port map (
            O => \N__48361\,
            I => \N__48350\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__48358\,
            I => \N__48350\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__48355\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__11317\ : Odrv4
    port map (
            O => \N__48350\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48345\,
            I => \N__48342\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__48342\,
            I => \N__48339\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__48339\,
            I => \N__48335\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48332\
        );

    \I__11312\ : Odrv4
    port map (
            O => \N__48335\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__48332\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__11310\ : CascadeMux
    port map (
            O => \N__48327\,
            I => \N__48324\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48321\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__48321\,
            I => \N__48318\
        );

    \I__11307\ : Span12Mux_v
    port map (
            O => \N__48318\,
            I => \N__48315\
        );

    \I__11306\ : Odrv12
    port map (
            O => \N__48315\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48312\,
            I => \N__48309\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48309\,
            I => \N__48304\
        );

    \I__11303\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48301\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48307\,
            I => \N__48298\
        );

    \I__11301\ : Span4Mux_v
    port map (
            O => \N__48304\,
            I => \N__48295\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48301\,
            I => \N__48292\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__48298\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__11298\ : Odrv4
    port map (
            O => \N__48295\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__11297\ : Odrv12
    port map (
            O => \N__48292\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48279\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48276\
        );

    \I__11294\ : InMux
    port map (
            O => \N__48283\,
            I => \N__48273\
        );

    \I__11293\ : InMux
    port map (
            O => \N__48282\,
            I => \N__48270\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__48279\,
            I => \N__48267\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__48276\,
            I => \N__48264\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__48273\,
            I => \N__48261\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__48270\,
            I => \N__48258\
        );

    \I__11288\ : Span4Mux_v
    port map (
            O => \N__48267\,
            I => \N__48249\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__48264\,
            I => \N__48249\
        );

    \I__11286\ : Span4Mux_v
    port map (
            O => \N__48261\,
            I => \N__48249\
        );

    \I__11285\ : Span4Mux_v
    port map (
            O => \N__48258\,
            I => \N__48249\
        );

    \I__11284\ : Odrv4
    port map (
            O => \N__48249\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__11283\ : CascadeMux
    port map (
            O => \N__48246\,
            I => \N__48243\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48240\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__48240\,
            I => \N__48237\
        );

    \I__11280\ : Span4Mux_v
    port map (
            O => \N__48237\,
            I => \N__48234\
        );

    \I__11279\ : Odrv4
    port map (
            O => \N__48234\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48231\,
            I => \N__48228\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__48228\,
            I => \N__48225\
        );

    \I__11276\ : Span4Mux_h
    port map (
            O => \N__48225\,
            I => \N__48222\
        );

    \I__11275\ : Span4Mux_v
    port map (
            O => \N__48222\,
            I => \N__48219\
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__48219\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48210\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48207\
        );

    \I__11271\ : CascadeMux
    port map (
            O => \N__48214\,
            I => \N__48204\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48201\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__48210\,
            I => \N__48196\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__48207\,
            I => \N__48196\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48204\,
            I => \N__48193\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__48201\,
            I => \N__48190\
        );

    \I__11265\ : Span4Mux_v
    port map (
            O => \N__48196\,
            I => \N__48185\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__48193\,
            I => \N__48185\
        );

    \I__11263\ : Span4Mux_h
    port map (
            O => \N__48190\,
            I => \N__48182\
        );

    \I__11262\ : Odrv4
    port map (
            O => \N__48185\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11261\ : Odrv4
    port map (
            O => \N__48182\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48174\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48174\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48167\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48164\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48167\,
            I => \N__48159\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__48164\,
            I => \N__48156\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48153\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48150\
        );

    \I__11252\ : Span4Mux_v
    port map (
            O => \N__48159\,
            I => \N__48143\
        );

    \I__11251\ : Span4Mux_v
    port map (
            O => \N__48156\,
            I => \N__48143\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__48153\,
            I => \N__48143\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48150\,
            I => \N__48140\
        );

    \I__11248\ : Span4Mux_h
    port map (
            O => \N__48143\,
            I => \N__48137\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__48140\,
            I => \N__48134\
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__48137\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__11245\ : Odrv4
    port map (
            O => \N__48134\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__11244\ : CascadeMux
    port map (
            O => \N__48129\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__11243\ : InMux
    port map (
            O => \N__48126\,
            I => \N__48123\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__48123\,
            I => \N__48120\
        );

    \I__11241\ : Odrv12
    port map (
            O => \N__48120\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48117\,
            I => \N__48113\
        );

    \I__11239\ : CascadeMux
    port map (
            O => \N__48116\,
            I => \N__48110\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48106\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48110\,
            I => \N__48103\
        );

    \I__11236\ : InMux
    port map (
            O => \N__48109\,
            I => \N__48100\
        );

    \I__11235\ : Odrv4
    port map (
            O => \N__48106\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__48103\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__48100\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__11232\ : CEMux
    port map (
            O => \N__48093\,
            I => \N__48090\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48090\,
            I => \N__48084\
        );

    \I__11230\ : CEMux
    port map (
            O => \N__48089\,
            I => \N__48081\
        );

    \I__11229\ : CEMux
    port map (
            O => \N__48088\,
            I => \N__48078\
        );

    \I__11228\ : CEMux
    port map (
            O => \N__48087\,
            I => \N__48075\
        );

    \I__11227\ : Span4Mux_h
    port map (
            O => \N__48084\,
            I => \N__48069\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48069\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48078\,
            I => \N__48066\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__48075\,
            I => \N__48063\
        );

    \I__11223\ : CEMux
    port map (
            O => \N__48074\,
            I => \N__48060\
        );

    \I__11222\ : Span4Mux_h
    port map (
            O => \N__48069\,
            I => \N__48057\
        );

    \I__11221\ : Span4Mux_v
    port map (
            O => \N__48066\,
            I => \N__48054\
        );

    \I__11220\ : Span4Mux_h
    port map (
            O => \N__48063\,
            I => \N__48051\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__48048\
        );

    \I__11218\ : Odrv4
    port map (
            O => \N__48057\,
            I => \delay_measurement_inst.delay_hc_timer.N_341_i\
        );

    \I__11217\ : Odrv4
    port map (
            O => \N__48054\,
            I => \delay_measurement_inst.delay_hc_timer.N_341_i\
        );

    \I__11216\ : Odrv4
    port map (
            O => \N__48051\,
            I => \delay_measurement_inst.delay_hc_timer.N_341_i\
        );

    \I__11215\ : Odrv4
    port map (
            O => \N__48048\,
            I => \delay_measurement_inst.delay_hc_timer.N_341_i\
        );

    \I__11214\ : InMux
    port map (
            O => \N__48039\,
            I => \N__48033\
        );

    \I__11213\ : InMux
    port map (
            O => \N__48038\,
            I => \N__48030\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48037\,
            I => \N__48027\
        );

    \I__11211\ : InMux
    port map (
            O => \N__48036\,
            I => \N__48024\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__48033\,
            I => \N__48019\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__48030\,
            I => \N__48019\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__48027\,
            I => \N__48016\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48024\,
            I => \N__48013\
        );

    \I__11206\ : Span4Mux_v
    port map (
            O => \N__48019\,
            I => \N__48010\
        );

    \I__11205\ : Odrv4
    port map (
            O => \N__48016\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__11204\ : Odrv12
    port map (
            O => \N__48013\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__11203\ : Odrv4
    port map (
            O => \N__48010\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__11202\ : InMux
    port map (
            O => \N__48003\,
            I => \N__48000\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__48000\,
            I => \N__47996\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47999\,
            I => \N__47993\
        );

    \I__11199\ : Span4Mux_h
    port map (
            O => \N__47996\,
            I => \N__47989\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47993\,
            I => \N__47986\
        );

    \I__11197\ : InMux
    port map (
            O => \N__47992\,
            I => \N__47983\
        );

    \I__11196\ : Span4Mux_v
    port map (
            O => \N__47989\,
            I => \N__47978\
        );

    \I__11195\ : Span4Mux_h
    port map (
            O => \N__47986\,
            I => \N__47978\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__47983\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__11193\ : Odrv4
    port map (
            O => \N__47978\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__11192\ : CascadeMux
    port map (
            O => \N__47973\,
            I => \N__47970\
        );

    \I__11191\ : InMux
    port map (
            O => \N__47970\,
            I => \N__47964\
        );

    \I__11190\ : InMux
    port map (
            O => \N__47969\,
            I => \N__47964\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__47964\,
            I => \N__47961\
        );

    \I__11188\ : Span4Mux_h
    port map (
            O => \N__47961\,
            I => \N__47958\
        );

    \I__11187\ : Odrv4
    port map (
            O => \N__47958\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__11186\ : CascadeMux
    port map (
            O => \N__47955\,
            I => \N__47951\
        );

    \I__11185\ : CascadeMux
    port map (
            O => \N__47954\,
            I => \N__47948\
        );

    \I__11184\ : InMux
    port map (
            O => \N__47951\,
            I => \N__47943\
        );

    \I__11183\ : InMux
    port map (
            O => \N__47948\,
            I => \N__47943\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47943\,
            I => \N__47940\
        );

    \I__11181\ : Span4Mux_v
    port map (
            O => \N__47940\,
            I => \N__47937\
        );

    \I__11180\ : Span4Mux_h
    port map (
            O => \N__47937\,
            I => \N__47934\
        );

    \I__11179\ : Odrv4
    port map (
            O => \N__47934\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__11178\ : InMux
    port map (
            O => \N__47931\,
            I => \N__47928\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__47928\,
            I => \N__47925\
        );

    \I__11176\ : Odrv12
    port map (
            O => \N__47925\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__11175\ : CascadeMux
    port map (
            O => \N__47922\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\
        );

    \I__11174\ : CascadeMux
    port map (
            O => \N__47919\,
            I => \N__47916\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47916\,
            I => \N__47913\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__47913\,
            I => \N__47910\
        );

    \I__11171\ : Odrv12
    port map (
            O => \N__47910\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47907\,
            I => \N__47904\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__47904\,
            I => \N__47901\
        );

    \I__11168\ : Span4Mux_h
    port map (
            O => \N__47901\,
            I => \N__47898\
        );

    \I__11167\ : Odrv4
    port map (
            O => \N__47898\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__11166\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47889\
        );

    \I__11165\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47889\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__47889\,
            I => \N__47884\
        );

    \I__11163\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47881\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47878\
        );

    \I__11161\ : Span4Mux_v
    port map (
            O => \N__47884\,
            I => \N__47875\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47881\,
            I => \N__47872\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__47878\,
            I => \N__47869\
        );

    \I__11158\ : Span4Mux_v
    port map (
            O => \N__47875\,
            I => \N__47866\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__47872\,
            I => \N__47861\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__47869\,
            I => \N__47861\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47866\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__47861\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__11153\ : InMux
    port map (
            O => \N__47856\,
            I => \N__47850\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47855\,
            I => \N__47847\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47854\,
            I => \N__47844\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47853\,
            I => \N__47841\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47850\,
            I => \N__47836\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47836\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47844\,
            I => \N__47833\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47841\,
            I => \N__47830\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__47836\,
            I => \N__47825\
        );

    \I__11144\ : Span4Mux_h
    port map (
            O => \N__47833\,
            I => \N__47825\
        );

    \I__11143\ : Odrv4
    port map (
            O => \N__47830\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__11142\ : Odrv4
    port map (
            O => \N__47825\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__11141\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47814\
        );

    \I__11140\ : InMux
    port map (
            O => \N__47819\,
            I => \N__47811\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47818\,
            I => \N__47808\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47817\,
            I => \N__47805\
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__47814\,
            I => \N__47802\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__47811\,
            I => \N__47799\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__47808\,
            I => \N__47794\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47794\
        );

    \I__11133\ : Span4Mux_h
    port map (
            O => \N__47802\,
            I => \N__47789\
        );

    \I__11132\ : Span4Mux_h
    port map (
            O => \N__47799\,
            I => \N__47789\
        );

    \I__11131\ : Odrv4
    port map (
            O => \N__47794\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11130\ : Odrv4
    port map (
            O => \N__47789\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__11129\ : CascadeMux
    port map (
            O => \N__47784\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__11128\ : CascadeMux
    port map (
            O => \N__47781\,
            I => \N__47778\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47775\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__47775\,
            I => \N__47772\
        );

    \I__11125\ : Span4Mux_h
    port map (
            O => \N__47772\,
            I => \N__47769\
        );

    \I__11124\ : Odrv4
    port map (
            O => \N__47769\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47763\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47760\
        );

    \I__11121\ : Sp12to4
    port map (
            O => \N__47760\,
            I => \N__47757\
        );

    \I__11120\ : Span12Mux_v
    port map (
            O => \N__47757\,
            I => \N__47754\
        );

    \I__11119\ : Span12Mux_h
    port map (
            O => \N__47754\,
            I => \N__47751\
        );

    \I__11118\ : Odrv12
    port map (
            O => \N__47751\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__11117\ : CascadeMux
    port map (
            O => \N__47748\,
            I => \N__47745\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47742\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__47742\,
            I => \N__47739\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__47739\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47736\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__11112\ : CascadeMux
    port map (
            O => \N__47733\,
            I => \N__47730\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47727\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__47727\,
            I => \N__47724\
        );

    \I__11109\ : Span12Mux_s7_h
    port map (
            O => \N__47724\,
            I => \N__47721\
        );

    \I__11108\ : Span12Mux_v
    port map (
            O => \N__47721\,
            I => \N__47718\
        );

    \I__11107\ : Span12Mux_h
    port map (
            O => \N__47718\,
            I => \N__47715\
        );

    \I__11106\ : Odrv12
    port map (
            O => \N__47715\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__11105\ : CascadeMux
    port map (
            O => \N__47712\,
            I => \N__47709\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47709\,
            I => \N__47706\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__47706\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47703\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47697\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47694\
        );

    \I__11099\ : Sp12to4
    port map (
            O => \N__47694\,
            I => \N__47691\
        );

    \I__11098\ : Span12Mux_h
    port map (
            O => \N__47691\,
            I => \N__47688\
        );

    \I__11097\ : Span12Mux_v
    port map (
            O => \N__47688\,
            I => \N__47685\
        );

    \I__11096\ : Odrv12
    port map (
            O => \N__47685\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47679\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47679\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47676\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__47673\,
            I => \N__47670\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47670\,
            I => \N__47667\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47667\,
            I => \N__47664\
        );

    \I__11089\ : Sp12to4
    port map (
            O => \N__47664\,
            I => \N__47661\
        );

    \I__11088\ : Span12Mux_h
    port map (
            O => \N__47661\,
            I => \N__47658\
        );

    \I__11087\ : Span12Mux_v
    port map (
            O => \N__47658\,
            I => \N__47655\
        );

    \I__11086\ : Odrv12
    port map (
            O => \N__47655\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__11085\ : CascadeMux
    port map (
            O => \N__47652\,
            I => \N__47649\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47649\,
            I => \N__47646\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__47646\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47643\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47637\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47634\
        );

    \I__11079\ : Span12Mux_h
    port map (
            O => \N__47634\,
            I => \N__47631\
        );

    \I__11078\ : Span12Mux_v
    port map (
            O => \N__47631\,
            I => \N__47628\
        );

    \I__11077\ : Odrv12
    port map (
            O => \N__47628\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__11076\ : CascadeMux
    port map (
            O => \N__47625\,
            I => \N__47622\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47619\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47619\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47616\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__11072\ : CascadeMux
    port map (
            O => \N__47613\,
            I => \N__47603\
        );

    \I__11071\ : CascadeMux
    port map (
            O => \N__47612\,
            I => \N__47599\
        );

    \I__11070\ : CascadeMux
    port map (
            O => \N__47611\,
            I => \N__47595\
        );

    \I__11069\ : CascadeMux
    port map (
            O => \N__47610\,
            I => \N__47591\
        );

    \I__11068\ : CascadeMux
    port map (
            O => \N__47609\,
            I => \N__47587\
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__47608\,
            I => \N__47584\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47607\,
            I => \N__47581\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47606\,
            I => \N__47566\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47603\,
            I => \N__47566\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47602\,
            I => \N__47566\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47599\,
            I => \N__47566\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47566\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47566\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47566\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47591\,
            I => \N__47563\
        );

    \I__11057\ : InMux
    port map (
            O => \N__47590\,
            I => \N__47556\
        );

    \I__11056\ : InMux
    port map (
            O => \N__47587\,
            I => \N__47556\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47584\,
            I => \N__47556\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47581\,
            I => \N__47553\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__47566\,
            I => \N__47546\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__47563\,
            I => \N__47546\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__47556\,
            I => \N__47546\
        );

    \I__11050\ : Span12Mux_h
    port map (
            O => \N__47553\,
            I => \N__47543\
        );

    \I__11049\ : Span12Mux_v
    port map (
            O => \N__47546\,
            I => \N__47540\
        );

    \I__11048\ : Odrv12
    port map (
            O => \N__47543\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__11047\ : Odrv12
    port map (
            O => \N__47540\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__11046\ : CascadeMux
    port map (
            O => \N__47535\,
            I => \N__47532\
        );

    \I__11045\ : InMux
    port map (
            O => \N__47532\,
            I => \N__47529\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__47529\,
            I => \N__47526\
        );

    \I__11043\ : Sp12to4
    port map (
            O => \N__47526\,
            I => \N__47523\
        );

    \I__11042\ : Span12Mux_h
    port map (
            O => \N__47523\,
            I => \N__47520\
        );

    \I__11041\ : Span12Mux_v
    port map (
            O => \N__47520\,
            I => \N__47517\
        );

    \I__11040\ : Odrv12
    port map (
            O => \N__47517\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__11039\ : CascadeMux
    port map (
            O => \N__47514\,
            I => \N__47511\
        );

    \I__11038\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47508\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__47508\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__11036\ : InMux
    port map (
            O => \N__47505\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47502\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__47496\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__11032\ : IoInMux
    port map (
            O => \N__47493\,
            I => \N__47490\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47490\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47487\,
            I => \N__47484\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__47484\,
            I => \N__47481\
        );

    \I__11028\ : Sp12to4
    port map (
            O => \N__47481\,
            I => \N__47478\
        );

    \I__11027\ : Span12Mux_v
    port map (
            O => \N__47478\,
            I => \N__47475\
        );

    \I__11026\ : Span12Mux_h
    port map (
            O => \N__47475\,
            I => \N__47472\
        );

    \I__11025\ : Odrv12
    port map (
            O => \N__47472\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__11024\ : CascadeMux
    port map (
            O => \N__47469\,
            I => \N__47466\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47466\,
            I => \N__47463\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47460\
        );

    \I__11021\ : Span4Mux_h
    port map (
            O => \N__47460\,
            I => \N__47457\
        );

    \I__11020\ : Span4Mux_h
    port map (
            O => \N__47457\,
            I => \N__47454\
        );

    \I__11019\ : Odrv4
    port map (
            O => \N__47454\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__11018\ : CascadeMux
    port map (
            O => \N__47451\,
            I => \N__47448\
        );

    \I__11017\ : InMux
    port map (
            O => \N__47448\,
            I => \N__47445\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__47445\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47442\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47439\,
            I => \N__47436\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__47436\,
            I => \N__47433\
        );

    \I__11012\ : Span12Mux_v
    port map (
            O => \N__47433\,
            I => \N__47430\
        );

    \I__11011\ : Span12Mux_h
    port map (
            O => \N__47430\,
            I => \N__47427\
        );

    \I__11010\ : Odrv12
    port map (
            O => \N__47427\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__11009\ : CascadeMux
    port map (
            O => \N__47424\,
            I => \N__47421\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47418\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__47418\,
            I => \N__47415\
        );

    \I__11006\ : Span4Mux_h
    port map (
            O => \N__47415\,
            I => \N__47412\
        );

    \I__11005\ : Span4Mux_h
    port map (
            O => \N__47412\,
            I => \N__47409\
        );

    \I__11004\ : Odrv4
    port map (
            O => \N__47409\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__47406\,
            I => \N__47403\
        );

    \I__11002\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47400\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__47400\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47397\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47391\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__47391\,
            I => \N__47388\
        );

    \I__10997\ : Span12Mux_s8_h
    port map (
            O => \N__47388\,
            I => \N__47385\
        );

    \I__10996\ : Span12Mux_h
    port map (
            O => \N__47385\,
            I => \N__47382\
        );

    \I__10995\ : Span12Mux_v
    port map (
            O => \N__47382\,
            I => \N__47379\
        );

    \I__10994\ : Odrv12
    port map (
            O => \N__47379\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__10993\ : CascadeMux
    port map (
            O => \N__47376\,
            I => \N__47373\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47373\,
            I => \N__47370\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__47370\,
            I => \N__47367\
        );

    \I__10990\ : Span4Mux_h
    port map (
            O => \N__47367\,
            I => \N__47364\
        );

    \I__10989\ : Span4Mux_h
    port map (
            O => \N__47364\,
            I => \N__47361\
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__47361\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__10987\ : CascadeMux
    port map (
            O => \N__47358\,
            I => \N__47355\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47355\,
            I => \N__47352\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47352\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__10984\ : InMux
    port map (
            O => \N__47349\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__10983\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47343\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__47343\,
            I => \N__47340\
        );

    \I__10981\ : Span12Mux_s9_h
    port map (
            O => \N__47340\,
            I => \N__47337\
        );

    \I__10980\ : Span12Mux_v
    port map (
            O => \N__47337\,
            I => \N__47334\
        );

    \I__10979\ : Span12Mux_h
    port map (
            O => \N__47334\,
            I => \N__47331\
        );

    \I__10978\ : Odrv12
    port map (
            O => \N__47331\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__10977\ : CascadeMux
    port map (
            O => \N__47328\,
            I => \N__47325\
        );

    \I__10976\ : InMux
    port map (
            O => \N__47325\,
            I => \N__47322\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47319\
        );

    \I__10974\ : Odrv4
    port map (
            O => \N__47319\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__10973\ : InMux
    port map (
            O => \N__47316\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47310\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__47310\,
            I => \N__47307\
        );

    \I__10970\ : Span12Mux_h
    port map (
            O => \N__47307\,
            I => \N__47304\
        );

    \I__10969\ : Span12Mux_v
    port map (
            O => \N__47304\,
            I => \N__47301\
        );

    \I__10968\ : Odrv12
    port map (
            O => \N__47301\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__10967\ : CascadeMux
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__10966\ : InMux
    port map (
            O => \N__47295\,
            I => \N__47292\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47292\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47289\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47286\,
            I => \N__47283\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47283\,
            I => \N__47280\
        );

    \I__10961\ : Span12Mux_h
    port map (
            O => \N__47280\,
            I => \N__47277\
        );

    \I__10960\ : Span12Mux_v
    port map (
            O => \N__47277\,
            I => \N__47274\
        );

    \I__10959\ : Odrv12
    port map (
            O => \N__47274\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__10958\ : CascadeMux
    port map (
            O => \N__47271\,
            I => \N__47268\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47265\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__47265\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47262\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__10954\ : CascadeMux
    port map (
            O => \N__47259\,
            I => \N__47256\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47253\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__47253\,
            I => \N__47250\
        );

    \I__10951\ : Span12Mux_h
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10950\ : Span12Mux_v
    port map (
            O => \N__47247\,
            I => \N__47244\
        );

    \I__10949\ : Odrv12
    port map (
            O => \N__47244\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__10948\ : CascadeMux
    port map (
            O => \N__47241\,
            I => \N__47238\
        );

    \I__10947\ : InMux
    port map (
            O => \N__47238\,
            I => \N__47235\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__47235\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47232\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__10944\ : CascadeMux
    port map (
            O => \N__47229\,
            I => \N__47226\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47223\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47223\,
            I => \N__47220\
        );

    \I__10941\ : Span12Mux_h
    port map (
            O => \N__47220\,
            I => \N__47217\
        );

    \I__10940\ : Span12Mux_v
    port map (
            O => \N__47217\,
            I => \N__47214\
        );

    \I__10939\ : Odrv12
    port map (
            O => \N__47214\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__47211\,
            I => \N__47208\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47208\,
            I => \N__47205\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__47205\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47202\,
            I => \bfn_18_23_0_\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47196\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__10932\ : CascadeMux
    port map (
            O => \N__47193\,
            I => \N__47190\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47187\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__47187\,
            I => \N__47184\
        );

    \I__10929\ : Odrv4
    port map (
            O => \N__47184\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47181\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_0_30\
        );

    \I__10927\ : CascadeMux
    port map (
            O => \N__47178\,
            I => \N__47175\
        );

    \I__10926\ : InMux
    port map (
            O => \N__47175\,
            I => \N__47169\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47169\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__47169\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO\
        );

    \I__10923\ : IoInMux
    port map (
            O => \N__47166\,
            I => \N__47137\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47124\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47124\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47124\
        );

    \I__10919\ : InMux
    port map (
            O => \N__47162\,
            I => \N__47124\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47161\,
            I => \N__47117\
        );

    \I__10917\ : InMux
    port map (
            O => \N__47160\,
            I => \N__47117\
        );

    \I__10916\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47117\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47108\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47108\
        );

    \I__10913\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47108\
        );

    \I__10912\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47108\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47098\
        );

    \I__10910\ : InMux
    port map (
            O => \N__47153\,
            I => \N__47098\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47098\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47098\
        );

    \I__10907\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47089\
        );

    \I__10906\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47089\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47089\
        );

    \I__10904\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47089\
        );

    \I__10903\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47082\
        );

    \I__10902\ : InMux
    port map (
            O => \N__47145\,
            I => \N__47082\
        );

    \I__10901\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47082\
        );

    \I__10900\ : InMux
    port map (
            O => \N__47143\,
            I => \N__47073\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47073\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47073\
        );

    \I__10897\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47073\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47070\
        );

    \I__10895\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47061\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47061\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47061\
        );

    \I__10892\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47061\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__47124\,
            I => \N__47056\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__47117\,
            I => \N__47056\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__47108\,
            I => \N__47053\
        );

    \I__10888\ : InMux
    port map (
            O => \N__47107\,
            I => \N__47050\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__47098\,
            I => \N__47047\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47040\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__47082\,
            I => \N__47040\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__47073\,
            I => \N__47040\
        );

    \I__10883\ : Span4Mux_s1_v
    port map (
            O => \N__47070\,
            I => \N__47037\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__47061\,
            I => \N__47034\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__47056\,
            I => \N__47029\
        );

    \I__10880\ : Span4Mux_v
    port map (
            O => \N__47053\,
            I => \N__47029\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47050\,
            I => \N__47022\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__47047\,
            I => \N__47022\
        );

    \I__10877\ : Span4Mux_v
    port map (
            O => \N__47040\,
            I => \N__47022\
        );

    \I__10876\ : Span4Mux_h
    port map (
            O => \N__47037\,
            I => \N__47019\
        );

    \I__10875\ : Span4Mux_h
    port map (
            O => \N__47034\,
            I => \N__47016\
        );

    \I__10874\ : Span4Mux_v
    port map (
            O => \N__47029\,
            I => \N__47011\
        );

    \I__10873\ : Span4Mux_v
    port map (
            O => \N__47022\,
            I => \N__47011\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__47019\,
            I => \N__47008\
        );

    \I__10871\ : Span4Mux_v
    port map (
            O => \N__47016\,
            I => \N__47005\
        );

    \I__10870\ : Span4Mux_h
    port map (
            O => \N__47011\,
            I => \N__47000\
        );

    \I__10869\ : Span4Mux_v
    port map (
            O => \N__47008\,
            I => \N__47000\
        );

    \I__10868\ : Odrv4
    port map (
            O => \N__47005\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__47000\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46995\,
            I => \N__46991\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46994\,
            I => \N__46988\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46991\,
            I => \N__46985\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46988\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30\
        );

    \I__10862\ : Odrv12
    port map (
            O => \N__46985\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46977\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46972\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46969\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46966\
        );

    \I__10857\ : Span4Mux_v
    port map (
            O => \N__46972\,
            I => \N__46961\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46969\,
            I => \N__46961\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46966\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10854\ : Odrv4
    port map (
            O => \N__46961\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46953\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46953\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46950\,
            I => \N__46947\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46947\,
            I => \N__46944\
        );

    \I__10849\ : Span4Mux_v
    port map (
            O => \N__46944\,
            I => \N__46940\
        );

    \I__10848\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46937\
        );

    \I__10847\ : Sp12to4
    port map (
            O => \N__46940\,
            I => \N__46933\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46929\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46926\
        );

    \I__10844\ : Span12Mux_h
    port map (
            O => \N__46933\,
            I => \N__46923\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46932\,
            I => \N__46920\
        );

    \I__10842\ : Span4Mux_v
    port map (
            O => \N__46929\,
            I => \N__46915\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46926\,
            I => \N__46915\
        );

    \I__10840\ : Odrv12
    port map (
            O => \N__46923\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46920\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__10838\ : Odrv4
    port map (
            O => \N__46915\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__10837\ : CascadeMux
    port map (
            O => \N__46908\,
            I => \N__46905\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46902\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__46902\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__10834\ : CascadeMux
    port map (
            O => \N__46899\,
            I => \N__46896\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46893\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46888\
        );

    \I__10831\ : CascadeMux
    port map (
            O => \N__46892\,
            I => \N__46885\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46882\
        );

    \I__10829\ : Span4Mux_v
    port map (
            O => \N__46888\,
            I => \N__46879\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46876\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46882\,
            I => \N__46873\
        );

    \I__10826\ : Sp12to4
    port map (
            O => \N__46879\,
            I => \N__46869\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__46876\,
            I => \N__46866\
        );

    \I__10824\ : Span4Mux_h
    port map (
            O => \N__46873\,
            I => \N__46863\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46860\
        );

    \I__10822\ : Span12Mux_h
    port map (
            O => \N__46869\,
            I => \N__46857\
        );

    \I__10821\ : Odrv4
    port map (
            O => \N__46866\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__10820\ : Odrv4
    port map (
            O => \N__46863\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46860\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__10818\ : Odrv12
    port map (
            O => \N__46857\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__10817\ : CascadeMux
    port map (
            O => \N__46848\,
            I => \N__46845\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46845\,
            I => \N__46842\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46842\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__10814\ : CascadeMux
    port map (
            O => \N__46839\,
            I => \N__46835\
        );

    \I__10813\ : CascadeMux
    port map (
            O => \N__46838\,
            I => \N__46832\
        );

    \I__10812\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46829\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46826\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46829\,
            I => \N__46822\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46826\,
            I => \N__46819\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46816\
        );

    \I__10807\ : Span4Mux_v
    port map (
            O => \N__46822\,
            I => \N__46813\
        );

    \I__10806\ : Span4Mux_v
    port map (
            O => \N__46819\,
            I => \N__46810\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46807\
        );

    \I__10804\ : Sp12to4
    port map (
            O => \N__46813\,
            I => \N__46801\
        );

    \I__10803\ : Sp12to4
    port map (
            O => \N__46810\,
            I => \N__46801\
        );

    \I__10802\ : Span4Mux_v
    port map (
            O => \N__46807\,
            I => \N__46798\
        );

    \I__10801\ : InMux
    port map (
            O => \N__46806\,
            I => \N__46795\
        );

    \I__10800\ : Span12Mux_h
    port map (
            O => \N__46801\,
            I => \N__46792\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__46798\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46795\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__10797\ : Odrv12
    port map (
            O => \N__46792\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__10796\ : CascadeMux
    port map (
            O => \N__46785\,
            I => \N__46771\
        );

    \I__10795\ : CascadeMux
    port map (
            O => \N__46784\,
            I => \N__46758\
        );

    \I__10794\ : CascadeMux
    port map (
            O => \N__46783\,
            I => \N__46755\
        );

    \I__10793\ : CascadeMux
    port map (
            O => \N__46782\,
            I => \N__46752\
        );

    \I__10792\ : CascadeMux
    port map (
            O => \N__46781\,
            I => \N__46745\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46742\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46729\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46778\,
            I => \N__46729\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46729\
        );

    \I__10787\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46729\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46729\
        );

    \I__10785\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46729\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46726\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46770\,
            I => \N__46721\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46769\,
            I => \N__46721\
        );

    \I__10781\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46714\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46714\
        );

    \I__10779\ : CascadeMux
    port map (
            O => \N__46766\,
            I => \N__46708\
        );

    \I__10778\ : CascadeMux
    port map (
            O => \N__46765\,
            I => \N__46705\
        );

    \I__10777\ : CascadeMux
    port map (
            O => \N__46764\,
            I => \N__46702\
        );

    \I__10776\ : InMux
    port map (
            O => \N__46763\,
            I => \N__46689\
        );

    \I__10775\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46689\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46689\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46758\,
            I => \N__46689\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46755\,
            I => \N__46689\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46752\,
            I => \N__46689\
        );

    \I__10770\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46686\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46683\
        );

    \I__10768\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46676\
        );

    \I__10767\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46676\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46676\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46673\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__46729\,
            I => \N__46668\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46726\,
            I => \N__46668\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46721\,
            I => \N__46665\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46720\,
            I => \N__46660\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46719\,
            I => \N__46660\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46657\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46644\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46644\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46711\,
            I => \N__46644\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46708\,
            I => \N__46644\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46705\,
            I => \N__46644\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46702\,
            I => \N__46644\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46689\,
            I => \N__46641\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__46686\,
            I => \N__46634\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46634\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__46676\,
            I => \N__46634\
        );

    \I__10748\ : Span4Mux_v
    port map (
            O => \N__46673\,
            I => \N__46629\
        );

    \I__10747\ : Span4Mux_v
    port map (
            O => \N__46668\,
            I => \N__46629\
        );

    \I__10746\ : Span12Mux_h
    port map (
            O => \N__46665\,
            I => \N__46624\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__46660\,
            I => \N__46624\
        );

    \I__10744\ : Span4Mux_h
    port map (
            O => \N__46657\,
            I => \N__46621\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46644\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10742\ : Odrv4
    port map (
            O => \N__46641\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__46634\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10740\ : Odrv4
    port map (
            O => \N__46629\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10739\ : Odrv12
    port map (
            O => \N__46624\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__46621\,
            I => \current_shift_inst.PI_CTRL.N_289\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46604\
        );

    \I__10736\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46601\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__46604\,
            I => \N__46598\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46601\,
            I => \N__46590\
        );

    \I__10733\ : Span4Mux_v
    port map (
            O => \N__46598\,
            I => \N__46586\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46597\,
            I => \N__46576\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46596\,
            I => \N__46571\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46595\,
            I => \N__46571\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46566\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46566\
        );

    \I__10727\ : Span4Mux_v
    port map (
            O => \N__46590\,
            I => \N__46557\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46553\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__46586\,
            I => \N__46550\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46547\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46525\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46525\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46582\,
            I => \N__46525\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46525\
        );

    \I__10719\ : InMux
    port map (
            O => \N__46580\,
            I => \N__46525\
        );

    \I__10718\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46525\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46576\,
            I => \N__46522\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46517\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__46566\,
            I => \N__46517\
        );

    \I__10714\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46503\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46503\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46503\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46503\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46561\,
            I => \N__46503\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46503\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__46557\,
            I => \N__46500\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46556\,
            I => \N__46497\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46553\,
            I => \N__46490\
        );

    \I__10705\ : Span4Mux_h
    port map (
            O => \N__46550\,
            I => \N__46490\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__46547\,
            I => \N__46490\
        );

    \I__10703\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46487\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46482\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46544\,
            I => \N__46482\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46543\,
            I => \N__46469\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46542\,
            I => \N__46469\
        );

    \I__10698\ : InMux
    port map (
            O => \N__46541\,
            I => \N__46469\
        );

    \I__10697\ : InMux
    port map (
            O => \N__46540\,
            I => \N__46469\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46539\,
            I => \N__46469\
        );

    \I__10695\ : InMux
    port map (
            O => \N__46538\,
            I => \N__46469\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__46525\,
            I => \N__46462\
        );

    \I__10693\ : Span4Mux_v
    port map (
            O => \N__46522\,
            I => \N__46462\
        );

    \I__10692\ : Span4Mux_v
    port map (
            O => \N__46517\,
            I => \N__46462\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46516\,
            I => \N__46459\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46452\
        );

    \I__10689\ : Span4Mux_h
    port map (
            O => \N__46500\,
            I => \N__46452\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__46497\,
            I => \N__46452\
        );

    \I__10687\ : Span4Mux_v
    port map (
            O => \N__46490\,
            I => \N__46449\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__46487\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__46482\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__46469\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10683\ : Odrv4
    port map (
            O => \N__46462\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46459\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__46452\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10680\ : Odrv4
    port map (
            O => \N__46449\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__10679\ : CascadeMux
    port map (
            O => \N__46434\,
            I => \N__46431\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46431\,
            I => \N__46428\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46428\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__10676\ : CascadeMux
    port map (
            O => \N__46425\,
            I => \N__46413\
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__46424\,
            I => \N__46410\
        );

    \I__10674\ : CascadeMux
    port map (
            O => \N__46423\,
            I => \N__46407\
        );

    \I__10673\ : CascadeMux
    port map (
            O => \N__46422\,
            I => \N__46404\
        );

    \I__10672\ : CascadeMux
    port map (
            O => \N__46421\,
            I => \N__46398\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46395\
        );

    \I__10670\ : CascadeMux
    port map (
            O => \N__46419\,
            I => \N__46380\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46375\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46359\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46359\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46359\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46359\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46359\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46404\,
            I => \N__46359\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46346\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46346\
        );

    \I__10660\ : InMux
    port map (
            O => \N__46401\,
            I => \N__46346\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46398\,
            I => \N__46346\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46395\,
            I => \N__46346\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46346\
        );

    \I__10656\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46343\
        );

    \I__10655\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46330\
        );

    \I__10654\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46330\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46330\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46330\
        );

    \I__10651\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46330\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46330\
        );

    \I__10649\ : CascadeMux
    port map (
            O => \N__46386\,
            I => \N__46326\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46323\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46320\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46315\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46315\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46312\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46309\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__46375\,
            I => \N__46306\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46374\,
            I => \N__46299\
        );

    \I__10640\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46299\
        );

    \I__10639\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46299\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46294\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46346\,
            I => \N__46294\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__46343\,
            I => \N__46289\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__46330\,
            I => \N__46289\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46329\,
            I => \N__46284\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46326\,
            I => \N__46284\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46323\,
            I => \N__46279\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__46320\,
            I => \N__46279\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__46315\,
            I => \N__46276\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46312\,
            I => \N__46263\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__46309\,
            I => \N__46263\
        );

    \I__10627\ : Span4Mux_v
    port map (
            O => \N__46306\,
            I => \N__46263\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__46299\,
            I => \N__46263\
        );

    \I__10625\ : Span4Mux_v
    port map (
            O => \N__46294\,
            I => \N__46263\
        );

    \I__10624\ : Span4Mux_v
    port map (
            O => \N__46289\,
            I => \N__46263\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__46284\,
            I => \N__46256\
        );

    \I__10622\ : Span12Mux_s10_v
    port map (
            O => \N__46279\,
            I => \N__46256\
        );

    \I__10621\ : Span12Mux_s7_h
    port map (
            O => \N__46276\,
            I => \N__46256\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__46263\,
            I => \N__46253\
        );

    \I__10619\ : Odrv12
    port map (
            O => \N__46256\,
            I => \current_shift_inst.PI_CTRL.N_290\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__46253\,
            I => \current_shift_inst.PI_CTRL.N_290\
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__46248\,
            I => \N__46245\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46245\,
            I => \N__46242\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__46242\,
            I => \N__46239\
        );

    \I__10614\ : Span4Mux_h
    port map (
            O => \N__46239\,
            I => \N__46236\
        );

    \I__10613\ : Span4Mux_v
    port map (
            O => \N__46236\,
            I => \N__46231\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46228\
        );

    \I__10611\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46225\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__46231\,
            I => \N__46220\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__46228\,
            I => \N__46220\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__46225\,
            I => \N__46214\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__46220\,
            I => \N__46214\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46211\
        );

    \I__10605\ : Span4Mux_h
    port map (
            O => \N__46214\,
            I => \N__46208\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__46211\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__10603\ : Odrv4
    port map (
            O => \N__46208\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46203\,
            I => \N__46200\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46200\,
            I => \N__46197\
        );

    \I__10600\ : Sp12to4
    port map (
            O => \N__46197\,
            I => \N__46194\
        );

    \I__10599\ : Span12Mux_h
    port map (
            O => \N__46194\,
            I => \N__46191\
        );

    \I__10598\ : Span12Mux_v
    port map (
            O => \N__46191\,
            I => \N__46188\
        );

    \I__10597\ : Odrv12
    port map (
            O => \N__46188\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__10596\ : CascadeMux
    port map (
            O => \N__46185\,
            I => \N__46182\
        );

    \I__10595\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__46179\,
            I => \N__46176\
        );

    \I__10593\ : Span4Mux_h
    port map (
            O => \N__46176\,
            I => \N__46173\
        );

    \I__10592\ : Span4Mux_h
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__46170\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__10590\ : CascadeMux
    port map (
            O => \N__46167\,
            I => \N__46164\
        );

    \I__10589\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46161\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__46161\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__46158\,
            I => \N__46155\
        );

    \I__10586\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46152\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__46152\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__10584\ : InMux
    port map (
            O => \N__46149\,
            I => \N__46146\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46143\
        );

    \I__10582\ : Span4Mux_v
    port map (
            O => \N__46143\,
            I => \N__46140\
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__46140\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__46137\,
            I => \N__46134\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46131\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__46131\,
            I => \N__46128\
        );

    \I__10577\ : Span4Mux_v
    port map (
            O => \N__46128\,
            I => \N__46125\
        );

    \I__10576\ : Odrv4
    port map (
            O => \N__46125\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46122\,
            I => \N__46119\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__46119\,
            I => \N__46116\
        );

    \I__10573\ : Odrv12
    port map (
            O => \N__46116\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__10572\ : CascadeMux
    port map (
            O => \N__46113\,
            I => \N__46110\
        );

    \I__10571\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46107\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__46107\,
            I => \N__46104\
        );

    \I__10569\ : Span4Mux_v
    port map (
            O => \N__46104\,
            I => \N__46101\
        );

    \I__10568\ : Odrv4
    port map (
            O => \N__46101\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46095\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__46095\,
            I => \N__46092\
        );

    \I__10565\ : Span4Mux_h
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__10564\ : Span4Mux_v
    port map (
            O => \N__46089\,
            I => \N__46086\
        );

    \I__10563\ : Odrv4
    port map (
            O => \N__46086\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__10562\ : CascadeMux
    port map (
            O => \N__46083\,
            I => \N__46080\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__46077\,
            I => \N__46074\
        );

    \I__10559\ : Span4Mux_h
    port map (
            O => \N__46074\,
            I => \N__46071\
        );

    \I__10558\ : Span4Mux_v
    port map (
            O => \N__46071\,
            I => \N__46068\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__46068\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__10556\ : InMux
    port map (
            O => \N__46065\,
            I => \N__46062\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46062\,
            I => \N__46059\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__46059\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__10553\ : CascadeMux
    port map (
            O => \N__46056\,
            I => \N__46053\
        );

    \I__10552\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46050\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46050\,
            I => \N__46047\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__46047\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__10549\ : InMux
    port map (
            O => \N__46044\,
            I => \N__46041\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__46041\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__46038\,
            I => \N__46035\
        );

    \I__10546\ : InMux
    port map (
            O => \N__46035\,
            I => \N__46032\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__46032\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46029\,
            I => \N__46026\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__46026\,
            I => \N__46023\
        );

    \I__10542\ : Span12Mux_h
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__10541\ : Odrv12
    port map (
            O => \N__46020\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__46017\,
            I => \N__46014\
        );

    \I__10539\ : InMux
    port map (
            O => \N__46014\,
            I => \N__46011\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46011\,
            I => \N__46008\
        );

    \I__10537\ : Span4Mux_h
    port map (
            O => \N__46008\,
            I => \N__46005\
        );

    \I__10536\ : Span4Mux_v
    port map (
            O => \N__46005\,
            I => \N__46002\
        );

    \I__10535\ : Span4Mux_v
    port map (
            O => \N__46002\,
            I => \N__45999\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__45999\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45992\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45989\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45992\,
            I => \N__45986\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__45989\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10529\ : Odrv4
    port map (
            O => \N__45986\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__45981\,
            I => \N__45978\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45975\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45975\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45969\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45969\,
            I => \N__45965\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45962\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__45965\,
            I => \N__45959\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__45962\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__45959\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45951\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45944\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45947\,
            I => \N__45941\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45944\,
            I => \N__45938\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__45941\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10513\ : Odrv4
    port map (
            O => \N__45938\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45930\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45930\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45924\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45920\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45917\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__45920\,
            I => \N__45914\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45917\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10505\ : Odrv4
    port map (
            O => \N__45914\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10504\ : CascadeMux
    port map (
            O => \N__45909\,
            I => \N__45906\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45903\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__45903\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45894\
        );

    \I__10499\ : Span4Mux_h
    port map (
            O => \N__45894\,
            I => \N__45891\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45891\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45888\,
            I => \N__45884\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45887\,
            I => \N__45881\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__45884\,
            I => \N__45878\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45881\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10493\ : Odrv4
    port map (
            O => \N__45878\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10492\ : CascadeMux
    port map (
            O => \N__45873\,
            I => \N__45870\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45867\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45867\,
            I => \N__45864\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__45864\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45857\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45854\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45857\,
            I => \N__45851\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45854\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__45851\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45846\,
            I => \N__45843\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45843\,
            I => \N__45840\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__45840\,
            I => \N__45837\
        );

    \I__10480\ : Span12Mux_v
    port map (
            O => \N__45837\,
            I => \N__45834\
        );

    \I__10479\ : Odrv12
    port map (
            O => \N__45834\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45828\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45828\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45825\,
            I => \N__45821\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45824\,
            I => \N__45818\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45821\,
            I => \N__45815\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45818\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10472\ : Odrv4
    port map (
            O => \N__45815\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__45807\,
            I => \N__45804\
        );

    \I__10469\ : Odrv12
    port map (
            O => \N__45804\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__10468\ : CascadeMux
    port map (
            O => \N__45801\,
            I => \N__45798\
        );

    \I__10467\ : InMux
    port map (
            O => \N__45798\,
            I => \N__45795\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45792\
        );

    \I__10465\ : Odrv4
    port map (
            O => \N__45792\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45789\,
            I => \N__45786\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__45786\,
            I => \N__45783\
        );

    \I__10462\ : Odrv12
    port map (
            O => \N__45783\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45780\,
            I => \N__45776\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45773\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45776\,
            I => \N__45770\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__45773\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10457\ : Odrv4
    port map (
            O => \N__45770\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45762\,
            I => \N__45759\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__10453\ : Odrv4
    port map (
            O => \N__45756\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45753\,
            I => \N__45750\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45746\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45743\
        );

    \I__10449\ : Span4Mux_v
    port map (
            O => \N__45746\,
            I => \N__45740\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__45743\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__45740\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__45735\,
            I => \N__45732\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__45729\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45723\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45723\,
            I => \N__45719\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45716\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__45719\,
            I => \N__45713\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45716\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__45713\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45705\
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__45705\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45699\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__45699\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45693\,
            I => \N__45689\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45686\
        );

    \I__10430\ : Span4Mux_v
    port map (
            O => \N__45689\,
            I => \N__45683\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45686\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10428\ : Odrv4
    port map (
            O => \N__45683\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10427\ : CascadeMux
    port map (
            O => \N__45678\,
            I => \N__45675\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45675\,
            I => \N__45672\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__45672\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45665\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45662\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45659\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__45662\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10420\ : Odrv4
    port map (
            O => \N__45659\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45651\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45651\,
            I => \N__45648\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__45648\,
            I => \N__45645\
        );

    \I__10416\ : Odrv4
    port map (
            O => \N__45645\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__10415\ : CascadeMux
    port map (
            O => \N__45642\,
            I => \N__45639\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45636\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__45636\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__45633\,
            I => \N__45630\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45627\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45624\
        );

    \I__10409\ : Span4Mux_h
    port map (
            O => \N__45624\,
            I => \N__45621\
        );

    \I__10408\ : Odrv4
    port map (
            O => \N__45621\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45618\,
            I => \N__45614\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45611\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__45614\,
            I => \N__45608\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45611\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10403\ : Odrv4
    port map (
            O => \N__45608\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45600\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45600\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__10400\ : CascadeMux
    port map (
            O => \N__45597\,
            I => \N__45594\
        );

    \I__10399\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45591\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45591\,
            I => \N__45588\
        );

    \I__10397\ : Span4Mux_v
    port map (
            O => \N__45588\,
            I => \N__45585\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__45585\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__10395\ : InMux
    port map (
            O => \N__45582\,
            I => \N__45578\
        );

    \I__10394\ : InMux
    port map (
            O => \N__45581\,
            I => \N__45575\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45572\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__45575\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10391\ : Odrv4
    port map (
            O => \N__45572\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10390\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45564\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45564\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__10388\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45558\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__45558\,
            I => \N__45554\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45551\
        );

    \I__10385\ : Odrv12
    port map (
            O => \N__45554\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45551\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10383\ : CascadeMux
    port map (
            O => \N__45546\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45537\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45532\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45532\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45529\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45537\,
            I => \N__45526\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__45532\,
            I => \N__45523\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45529\,
            I => \N__45520\
        );

    \I__10375\ : Odrv12
    port map (
            O => \N__45526\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45523\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__45520\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10372\ : CascadeMux
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45504\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45504\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__45504\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45497\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45494\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__45497\,
            I => \N__45490\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__45494\,
            I => \N__45487\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45484\
        );

    \I__10363\ : Span4Mux_h
    port map (
            O => \N__45490\,
            I => \N__45481\
        );

    \I__10362\ : Span4Mux_v
    port map (
            O => \N__45487\,
            I => \N__45478\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__45484\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__10360\ : Odrv4
    port map (
            O => \N__45481\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__10359\ : Odrv4
    port map (
            O => \N__45478\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__10358\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45467\
        );

    \I__10357\ : InMux
    port map (
            O => \N__45470\,
            I => \N__45463\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45467\,
            I => \N__45459\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45466\,
            I => \N__45456\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__45463\,
            I => \N__45453\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45450\
        );

    \I__10352\ : Span4Mux_v
    port map (
            O => \N__45459\,
            I => \N__45443\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__45456\,
            I => \N__45443\
        );

    \I__10350\ : Span4Mux_h
    port map (
            O => \N__45453\,
            I => \N__45443\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45450\,
            I => \N__45440\
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__45443\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__45440\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45429\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45429\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45429\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45419\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45419\
        );

    \I__10341\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45416\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__45419\,
            I => \N__45412\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__45416\,
            I => \N__45409\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45406\
        );

    \I__10337\ : Span4Mux_v
    port map (
            O => \N__45412\,
            I => \N__45403\
        );

    \I__10336\ : Span4Mux_v
    port map (
            O => \N__45409\,
            I => \N__45398\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__45406\,
            I => \N__45398\
        );

    \I__10334\ : Odrv4
    port map (
            O => \N__45403\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__45398\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45390\,
            I => \N__45387\
        );

    \I__10330\ : Span4Mux_h
    port map (
            O => \N__45387\,
            I => \N__45384\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__45384\,
            I => \N__45380\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45377\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__45380\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45377\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45369\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45369\,
            I => \N__45365\
        );

    \I__10323\ : InMux
    port map (
            O => \N__45368\,
            I => \N__45361\
        );

    \I__10322\ : Span4Mux_h
    port map (
            O => \N__45365\,
            I => \N__45358\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45355\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45361\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10319\ : Odrv4
    port map (
            O => \N__45358\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__45355\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45342\
        );

    \I__10316\ : InMux
    port map (
            O => \N__45347\,
            I => \N__45339\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45336\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45333\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45342\,
            I => \N__45330\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__45339\,
            I => \N__45327\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45336\,
            I => \N__45324\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__45333\,
            I => \N__45321\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__45330\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10308\ : Odrv4
    port map (
            O => \N__45327\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10307\ : Odrv4
    port map (
            O => \N__45324\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10306\ : Odrv4
    port map (
            O => \N__45321\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__45312\,
            I => \N__45307\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45311\,
            I => \N__45304\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45299\
        );

    \I__10302\ : InMux
    port map (
            O => \N__45307\,
            I => \N__45299\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__45304\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45299\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45289\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45293\,
            I => \N__45284\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45292\,
            I => \N__45284\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45289\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__45284\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45276\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__45276\,
            I => \N__45271\
        );

    \I__10292\ : InMux
    port map (
            O => \N__45275\,
            I => \N__45268\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45274\,
            I => \N__45265\
        );

    \I__10290\ : Span4Mux_v
    port map (
            O => \N__45271\,
            I => \N__45262\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45268\,
            I => \N__45259\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45265\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__45262\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10286\ : Odrv4
    port map (
            O => \N__45259\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45248\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45243\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__45248\,
            I => \N__45240\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45235\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45246\,
            I => \N__45235\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__45243\,
            I => \N__45232\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__45240\,
            I => \N__45227\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45227\
        );

    \I__10277\ : Odrv12
    port map (
            O => \N__45232\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__45227\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10275\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45216\
        );

    \I__10274\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45216\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__45216\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__10272\ : CascadeMux
    port map (
            O => \N__45213\,
            I => \N__45210\
        );

    \I__10271\ : InMux
    port map (
            O => \N__45210\,
            I => \N__45205\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45209\,
            I => \N__45202\
        );

    \I__10269\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45199\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__45205\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__45202\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45199\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10265\ : CascadeMux
    port map (
            O => \N__45192\,
            I => \N__45187\
        );

    \I__10264\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45184\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45180\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45177\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45174\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45183\,
            I => \N__45171\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__45180\,
            I => \N__45168\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45177\,
            I => \N__45165\
        );

    \I__10257\ : Span4Mux_h
    port map (
            O => \N__45174\,
            I => \N__45162\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45171\,
            I => \N__45159\
        );

    \I__10255\ : Span4Mux_v
    port map (
            O => \N__45168\,
            I => \N__45156\
        );

    \I__10254\ : Span4Mux_h
    port map (
            O => \N__45165\,
            I => \N__45153\
        );

    \I__10253\ : Span4Mux_v
    port map (
            O => \N__45162\,
            I => \N__45148\
        );

    \I__10252\ : Span4Mux_h
    port map (
            O => \N__45159\,
            I => \N__45148\
        );

    \I__10251\ : Odrv4
    port map (
            O => \N__45156\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10250\ : Odrv4
    port map (
            O => \N__45153\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__45148\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45141\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__10247\ : CascadeMux
    port map (
            O => \N__45138\,
            I => \N__45135\
        );

    \I__10246\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45130\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45127\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45124\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__45130\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__45127\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__45124\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45117\,
            I => \bfn_18_13_0_\
        );

    \I__10239\ : CascadeMux
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45111\,
            I => \N__45106\
        );

    \I__10237\ : InMux
    port map (
            O => \N__45110\,
            I => \N__45103\
        );

    \I__10236\ : InMux
    port map (
            O => \N__45109\,
            I => \N__45100\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45106\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__45103\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__45100\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10232\ : InMux
    port map (
            O => \N__45093\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__10231\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45086\
        );

    \I__10230\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45083\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__45086\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45083\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10227\ : CascadeMux
    port map (
            O => \N__45078\,
            I => \N__45075\
        );

    \I__10226\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45070\
        );

    \I__10225\ : InMux
    port map (
            O => \N__45074\,
            I => \N__45067\
        );

    \I__10224\ : InMux
    port map (
            O => \N__45073\,
            I => \N__45064\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__45070\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__45067\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__45064\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10220\ : InMux
    port map (
            O => \N__45057\,
            I => \N__45052\
        );

    \I__10219\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45049\
        );

    \I__10218\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45046\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45042\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__45049\,
            I => \N__45037\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__45046\,
            I => \N__45037\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45045\,
            I => \N__45034\
        );

    \I__10213\ : Span4Mux_h
    port map (
            O => \N__45042\,
            I => \N__45027\
        );

    \I__10212\ : Span4Mux_v
    port map (
            O => \N__45037\,
            I => \N__45027\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__45034\,
            I => \N__45027\
        );

    \I__10210\ : Span4Mux_h
    port map (
            O => \N__45027\,
            I => \N__45024\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__45024\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__10208\ : InMux
    port map (
            O => \N__45021\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__10207\ : InMux
    port map (
            O => \N__45018\,
            I => \N__45014\
        );

    \I__10206\ : InMux
    port map (
            O => \N__45017\,
            I => \N__45011\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__45014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__45011\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__45006\,
            I => \N__45003\
        );

    \I__10202\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44998\
        );

    \I__10201\ : InMux
    port map (
            O => \N__45002\,
            I => \N__44995\
        );

    \I__10200\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44992\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__44998\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__44995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44992\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44979\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44976\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44971\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44971\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44979\,
            I => \N__44968\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__44976\,
            I => \N__44965\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44971\,
            I => \N__44962\
        );

    \I__10189\ : Span4Mux_h
    port map (
            O => \N__44968\,
            I => \N__44959\
        );

    \I__10188\ : Span4Mux_v
    port map (
            O => \N__44965\,
            I => \N__44956\
        );

    \I__10187\ : Span4Mux_h
    port map (
            O => \N__44962\,
            I => \N__44953\
        );

    \I__10186\ : Odrv4
    port map (
            O => \N__44959\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__44956\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__44953\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44946\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44943\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44937\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44933\
        );

    \I__10179\ : CascadeMux
    port map (
            O => \N__44936\,
            I => \N__44930\
        );

    \I__10178\ : Span4Mux_v
    port map (
            O => \N__44933\,
            I => \N__44926\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44923\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44920\
        );

    \I__10175\ : Odrv4
    port map (
            O => \N__44926\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44923\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44920\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44908\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44912\,
            I => \N__44903\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44903\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44908\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44903\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10167\ : CascadeMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44888\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44888\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44885\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44888\,
            I => \N__44882\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44885\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10161\ : Odrv4
    port map (
            O => \N__44882\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10160\ : CascadeMux
    port map (
            O => \N__44877\,
            I => \N__44874\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44869\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44873\,
            I => \N__44866\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44863\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44869\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44866\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44863\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44856\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__44853\,
            I => \N__44850\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44845\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44842\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44839\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__44845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__44842\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44839\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44832\,
            I => \bfn_18_12_0_\
        );

    \I__10144\ : CascadeMux
    port map (
            O => \N__44829\,
            I => \N__44826\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44826\,
            I => \N__44821\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44825\,
            I => \N__44818\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44815\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44821\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44818\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10137\ : CascadeMux
    port map (
            O => \N__44808\,
            I => \N__44802\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44799\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44806\,
            I => \N__44796\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44793\
        );

    \I__10133\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44790\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44799\,
            I => \N__44781\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44781\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44793\,
            I => \N__44781\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44790\,
            I => \N__44781\
        );

    \I__10128\ : Span4Mux_v
    port map (
            O => \N__44781\,
            I => \N__44778\
        );

    \I__10127\ : Odrv4
    port map (
            O => \N__44778\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44775\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__10125\ : CascadeMux
    port map (
            O => \N__44772\,
            I => \N__44769\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44764\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44761\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44758\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44764\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__44761\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44758\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44751\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__10117\ : CascadeMux
    port map (
            O => \N__44748\,
            I => \N__44745\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44740\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44737\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44743\,
            I => \N__44734\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__44737\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__44734\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44727\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__10109\ : CascadeMux
    port map (
            O => \N__44724\,
            I => \N__44721\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44716\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44713\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44710\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__44716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__44713\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10102\ : InMux
    port map (
            O => \N__44703\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__10101\ : CascadeMux
    port map (
            O => \N__44700\,
            I => \N__44697\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44692\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44689\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44695\,
            I => \N__44686\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44692\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44689\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10094\ : InMux
    port map (
            O => \N__44679\,
            I => \N__44675\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44672\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44675\,
            I => \N__44665\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__44672\,
            I => \N__44665\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44671\,
            I => \N__44662\
        );

    \I__10089\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44659\
        );

    \I__10088\ : Span4Mux_v
    port map (
            O => \N__44665\,
            I => \N__44654\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44662\,
            I => \N__44654\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__44659\,
            I => \N__44651\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__44654\,
            I => \N__44648\
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__44651\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__44648\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44643\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__10081\ : CascadeMux
    port map (
            O => \N__44640\,
            I => \N__44637\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44637\,
            I => \N__44632\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44629\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44626\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44632\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__44629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44626\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10074\ : CascadeMux
    port map (
            O => \N__44619\,
            I => \N__44614\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44618\,
            I => \N__44610\
        );

    \I__10072\ : InMux
    port map (
            O => \N__44617\,
            I => \N__44607\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44614\,
            I => \N__44604\
        );

    \I__10070\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44601\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__44610\,
            I => \N__44596\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44607\,
            I => \N__44596\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__44604\,
            I => \N__44593\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__44601\,
            I => \N__44590\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__44596\,
            I => \N__44587\
        );

    \I__10064\ : Span4Mux_h
    port map (
            O => \N__44593\,
            I => \N__44584\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__44590\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10062\ : Odrv4
    port map (
            O => \N__44587\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__44584\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44577\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__10059\ : CascadeMux
    port map (
            O => \N__44574\,
            I => \N__44571\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44566\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44563\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44560\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__44566\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44563\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__44560\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44553\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__10051\ : CascadeMux
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44542\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44539\
        );

    \I__10048\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44536\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44542\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44539\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44536\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44529\,
            I => \bfn_18_11_0_\
        );

    \I__10043\ : CascadeMux
    port map (
            O => \N__44526\,
            I => \N__44523\
        );

    \I__10042\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44518\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44515\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44521\,
            I => \N__44512\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__44518\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44515\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__44512\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44505\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__10035\ : CascadeMux
    port map (
            O => \N__44502\,
            I => \N__44499\
        );

    \I__10034\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44494\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44491\
        );

    \I__10032\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44488\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44494\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44491\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__44488\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44481\,
            I => \N__44476\
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__44480\,
            I => \N__44472\
        );

    \I__10026\ : CascadeMux
    port map (
            O => \N__44479\,
            I => \N__44469\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__44476\,
            I => \N__44466\
        );

    \I__10024\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44459\
        );

    \I__10023\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44459\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44459\
        );

    \I__10021\ : Span4Mux_v
    port map (
            O => \N__44466\,
            I => \N__44456\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__44459\,
            I => \N__44453\
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__44456\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10018\ : Odrv4
    port map (
            O => \N__44453\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10017\ : InMux
    port map (
            O => \N__44448\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__10016\ : CascadeMux
    port map (
            O => \N__44445\,
            I => \N__44442\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44442\,
            I => \N__44437\
        );

    \I__10014\ : InMux
    port map (
            O => \N__44441\,
            I => \N__44434\
        );

    \I__10013\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44431\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44434\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__44431\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44424\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__44421\,
            I => \N__44418\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44413\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44410\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44416\,
            I => \N__44407\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44407\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44400\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__44397\,
            I => \N__44394\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44389\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44386\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44383\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__44389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__44386\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44383\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44376\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9992\ : CascadeMux
    port map (
            O => \N__44373\,
            I => \N__44370\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44370\,
            I => \N__44365\
        );

    \I__9990\ : InMux
    port map (
            O => \N__44369\,
            I => \N__44362\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44359\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44365\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__44362\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__44359\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44352\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9984\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44342\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44339\
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__44342\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__44339\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__9979\ : CascadeMux
    port map (
            O => \N__44334\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\
        );

    \I__9978\ : InMux
    port map (
            O => \N__44331\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9977\ : CascadeMux
    port map (
            O => \N__44328\,
            I => \N__44325\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44320\
        );

    \I__9975\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44317\
        );

    \I__9974\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44314\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44320\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__44317\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__44314\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44307\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9969\ : CascadeMux
    port map (
            O => \N__44304\,
            I => \N__44301\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44296\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44300\,
            I => \N__44293\
        );

    \I__9966\ : InMux
    port map (
            O => \N__44299\,
            I => \N__44290\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44296\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__44293\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44290\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9962\ : InMux
    port map (
            O => \N__44283\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9961\ : CascadeMux
    port map (
            O => \N__44280\,
            I => \N__44277\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44277\,
            I => \N__44272\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44269\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44266\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44272\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__44269\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44266\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44259\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9953\ : CascadeMux
    port map (
            O => \N__44256\,
            I => \N__44253\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44253\,
            I => \N__44248\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44245\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44251\,
            I => \N__44242\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__44248\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__44245\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__44242\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9946\ : InMux
    port map (
            O => \N__44235\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9945\ : CascadeMux
    port map (
            O => \N__44232\,
            I => \N__44229\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44229\,
            I => \N__44224\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44221\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44218\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__44224\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44221\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44218\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44211\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__44208\,
            I => \N__44205\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44200\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__44204\,
            I => \N__44197\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44194\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__44200\,
            I => \N__44191\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44188\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44194\,
            I => \N__44185\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__44191\,
            I => \N__44180\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44188\,
            I => \N__44180\
        );

    \I__9928\ : Span12Mux_s4_v
    port map (
            O => \N__44185\,
            I => \N__44177\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__44180\,
            I => \N__44174\
        );

    \I__9926\ : Odrv12
    port map (
            O => \N__44177\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__44174\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44165\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__44165\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__44162\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__44157\,
            I => \N__44154\
        );

    \I__9919\ : InMux
    port map (
            O => \N__44154\,
            I => \N__44151\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44151\,
            I => \N__44148\
        );

    \I__9917\ : Odrv12
    port map (
            O => \N__44148\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44145\,
            I => \N__44141\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__44144\,
            I => \N__44138\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__44141\,
            I => \N__44134\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44131\
        );

    \I__9912\ : CascadeMux
    port map (
            O => \N__44137\,
            I => \N__44128\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__44134\,
            I => \N__44121\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44131\,
            I => \N__44121\
        );

    \I__9909\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44118\
        );

    \I__9908\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44115\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44112\
        );

    \I__9906\ : Span4Mux_h
    port map (
            O => \N__44121\,
            I => \N__44107\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44118\,
            I => \N__44107\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__44115\,
            I => \N__44104\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__44112\,
            I => \N__44101\
        );

    \I__9902\ : Span4Mux_h
    port map (
            O => \N__44107\,
            I => \N__44098\
        );

    \I__9901\ : Span12Mux_h
    port map (
            O => \N__44104\,
            I => \N__44095\
        );

    \I__9900\ : Span12Mux_v
    port map (
            O => \N__44101\,
            I => \N__44092\
        );

    \I__9899\ : Span4Mux_v
    port map (
            O => \N__44098\,
            I => \N__44089\
        );

    \I__9898\ : Odrv12
    port map (
            O => \N__44095\,
            I => \phase_controller_inst2.start_latched\
        );

    \I__9897\ : Odrv12
    port map (
            O => \N__44092\,
            I => \phase_controller_inst2.start_latched\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__44089\,
            I => \phase_controller_inst2.start_latched\
        );

    \I__9895\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44078\
        );

    \I__9894\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44075\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__44078\,
            I => \N__44069\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44069\
        );

    \I__9891\ : InMux
    port map (
            O => \N__44074\,
            I => \N__44066\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__44069\,
            I => \N__44063\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__44066\,
            I => \phase_controller_inst2.running\
        );

    \I__9888\ : Odrv4
    port map (
            O => \N__44063\,
            I => \phase_controller_inst2.running\
        );

    \I__9887\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44052\
        );

    \I__9886\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44052\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44049\
        );

    \I__9884\ : Odrv12
    port map (
            O => \N__44049\,
            I => \phase_controller_inst2.N_39\
        );

    \I__9883\ : CEMux
    port map (
            O => \N__44046\,
            I => \N__44043\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__44040\
        );

    \I__9881\ : Odrv12
    port map (
            O => \N__44040\,
            I => \phase_controller_inst2.stoper_tr.N_39_0\
        );

    \I__9880\ : InMux
    port map (
            O => \N__44037\,
            I => \N__44031\
        );

    \I__9879\ : InMux
    port map (
            O => \N__44036\,
            I => \N__44031\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__44031\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__9877\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44025\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__44022\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__44022\,
            I => \N__44019\
        );

    \I__9874\ : Odrv4
    port map (
            O => \N__44019\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__9873\ : InMux
    port map (
            O => \N__44016\,
            I => \N__44013\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__44013\,
            I => \N__44010\
        );

    \I__9871\ : Span4Mux_v
    port map (
            O => \N__44010\,
            I => \N__44007\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__44007\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__9869\ : InMux
    port map (
            O => \N__44004\,
            I => \N__44001\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__44001\,
            I => \N__43998\
        );

    \I__9867\ : Span4Mux_h
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__9866\ : Odrv4
    port map (
            O => \N__43995\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__9865\ : CascadeMux
    port map (
            O => \N__43992\,
            I => \N__43989\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43989\,
            I => \N__43986\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43986\,
            I => \N__43983\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__43983\,
            I => \N__43980\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__43980\,
            I => \N__43974\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43971\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43978\,
            I => \N__43968\
        );

    \I__9858\ : CascadeMux
    port map (
            O => \N__43977\,
            I => \N__43965\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__43974\,
            I => \N__43962\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__43971\,
            I => \N__43957\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43968\,
            I => \N__43957\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43965\,
            I => \N__43954\
        );

    \I__9853\ : Span4Mux_h
    port map (
            O => \N__43962\,
            I => \N__43951\
        );

    \I__9852\ : Span4Mux_h
    port map (
            O => \N__43957\,
            I => \N__43948\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__43954\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9850\ : Odrv4
    port map (
            O => \N__43951\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__43948\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43941\,
            I => \N__43938\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43938\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43935\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__9845\ : CascadeMux
    port map (
            O => \N__43932\,
            I => \N__43929\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43926\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43926\,
            I => \N__43923\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__43923\,
            I => \N__43919\
        );

    \I__9841\ : CascadeMux
    port map (
            O => \N__43922\,
            I => \N__43916\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__43919\,
            I => \N__43912\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43909\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43906\
        );

    \I__9837\ : Span4Mux_h
    port map (
            O => \N__43912\,
            I => \N__43902\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43909\,
            I => \N__43897\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43906\,
            I => \N__43897\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43894\
        );

    \I__9833\ : Span4Mux_h
    port map (
            O => \N__43902\,
            I => \N__43891\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__43897\,
            I => \N__43888\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__43894\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9830\ : Odrv4
    port map (
            O => \N__43891\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9829\ : Odrv4
    port map (
            O => \N__43888\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43878\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43875\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__9825\ : CascadeMux
    port map (
            O => \N__43872\,
            I => \N__43869\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43862\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__43865\,
            I => \N__43859\
        );

    \I__9821\ : Span4Mux_v
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43852\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43849\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43846\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43852\,
            I => \N__43843\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__43849\,
            I => \N__43835\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43846\,
            I => \N__43835\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__43843\,
            I => \N__43835\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43842\,
            I => \N__43832\
        );

    \I__9812\ : Span4Mux_h
    port map (
            O => \N__43835\,
            I => \N__43829\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__43832\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__43829\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__43824\,
            I => \N__43821\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43818\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43818\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43815\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__9805\ : CascadeMux
    port map (
            O => \N__43812\,
            I => \N__43809\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43809\,
            I => \N__43806\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43806\,
            I => \N__43803\
        );

    \I__9802\ : Span4Mux_v
    port map (
            O => \N__43803\,
            I => \N__43798\
        );

    \I__9801\ : CascadeMux
    port map (
            O => \N__43802\,
            I => \N__43795\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43792\
        );

    \I__9799\ : Span4Mux_v
    port map (
            O => \N__43798\,
            I => \N__43789\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43795\,
            I => \N__43786\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__43792\,
            I => \N__43782\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__43789\,
            I => \N__43779\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43786\,
            I => \N__43776\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43785\,
            I => \N__43773\
        );

    \I__9793\ : Span4Mux_v
    port map (
            O => \N__43782\,
            I => \N__43770\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__43779\,
            I => \N__43765\
        );

    \I__9791\ : Span4Mux_v
    port map (
            O => \N__43776\,
            I => \N__43765\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43773\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__43770\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9788\ : Odrv4
    port map (
            O => \N__43765\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9787\ : CascadeMux
    port map (
            O => \N__43758\,
            I => \N__43755\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43755\,
            I => \N__43752\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__43752\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43749\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43746\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43740\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43740\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43737\,
            I => \N__43734\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43734\,
            I => \N__43731\
        );

    \I__9778\ : Span4Mux_h
    port map (
            O => \N__43731\,
            I => \N__43728\
        );

    \I__9777\ : Sp12to4
    port map (
            O => \N__43728\,
            I => \N__43725\
        );

    \I__9776\ : Span12Mux_v
    port map (
            O => \N__43725\,
            I => \N__43722\
        );

    \I__9775\ : Span12Mux_h
    port map (
            O => \N__43722\,
            I => \N__43719\
        );

    \I__9774\ : Odrv12
    port map (
            O => \N__43719\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__43716\,
            I => \N__43713\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43710\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43704\,
            I => \phase_controller_inst1.stateZ0Z_5\
        );

    \I__9768\ : IoInMux
    port map (
            O => \N__43701\,
            I => \N__43697\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43694\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__43697\,
            I => test_c
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43694\,
            I => test_c
        );

    \I__9764\ : InMux
    port map (
            O => \N__43689\,
            I => \N__43683\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43683\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43683\,
            I => \N__43680\
        );

    \I__9761\ : Span4Mux_s3_v
    port map (
            O => \N__43680\,
            I => \N__43677\
        );

    \I__9760\ : Span4Mux_h
    port map (
            O => \N__43677\,
            I => \N__43673\
        );

    \I__9759\ : CEMux
    port map (
            O => \N__43676\,
            I => \N__43670\
        );

    \I__9758\ : Span4Mux_h
    port map (
            O => \N__43673\,
            I => \N__43664\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43664\
        );

    \I__9756\ : CEMux
    port map (
            O => \N__43669\,
            I => \N__43660\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__43664\,
            I => \N__43656\
        );

    \I__9754\ : CEMux
    port map (
            O => \N__43663\,
            I => \N__43653\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43660\,
            I => \N__43650\
        );

    \I__9752\ : CEMux
    port map (
            O => \N__43659\,
            I => \N__43647\
        );

    \I__9751\ : Span4Mux_h
    port map (
            O => \N__43656\,
            I => \N__43642\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__43653\,
            I => \N__43642\
        );

    \I__9749\ : Span4Mux_s1_v
    port map (
            O => \N__43650\,
            I => \N__43638\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43635\
        );

    \I__9747\ : Span4Mux_v
    port map (
            O => \N__43642\,
            I => \N__43632\
        );

    \I__9746\ : CEMux
    port map (
            O => \N__43641\,
            I => \N__43629\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__43638\,
            I => \N__43620\
        );

    \I__9744\ : Span4Mux_h
    port map (
            O => \N__43635\,
            I => \N__43620\
        );

    \I__9743\ : Span4Mux_v
    port map (
            O => \N__43632\,
            I => \N__43617\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43629\,
            I => \N__43614\
        );

    \I__9741\ : CEMux
    port map (
            O => \N__43628\,
            I => \N__43611\
        );

    \I__9740\ : CEMux
    port map (
            O => \N__43627\,
            I => \N__43608\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43603\
        );

    \I__9738\ : CEMux
    port map (
            O => \N__43625\,
            I => \N__43600\
        );

    \I__9737\ : Sp12to4
    port map (
            O => \N__43620\,
            I => \N__43596\
        );

    \I__9736\ : Sp12to4
    port map (
            O => \N__43617\,
            I => \N__43591\
        );

    \I__9735\ : Sp12to4
    port map (
            O => \N__43614\,
            I => \N__43591\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43588\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43585\
        );

    \I__9732\ : CEMux
    port map (
            O => \N__43607\,
            I => \N__43582\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43579\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43603\,
            I => \N__43574\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43600\,
            I => \N__43574\
        );

    \I__9728\ : CEMux
    port map (
            O => \N__43599\,
            I => \N__43571\
        );

    \I__9727\ : Span12Mux_s11_v
    port map (
            O => \N__43596\,
            I => \N__43566\
        );

    \I__9726\ : Span12Mux_h
    port map (
            O => \N__43591\,
            I => \N__43566\
        );

    \I__9725\ : Span4Mux_h
    port map (
            O => \N__43588\,
            I => \N__43559\
        );

    \I__9724\ : Span4Mux_h
    port map (
            O => \N__43585\,
            I => \N__43559\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__43582\,
            I => \N__43559\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__43579\,
            I => \N__43556\
        );

    \I__9721\ : Span4Mux_h
    port map (
            O => \N__43574\,
            I => \N__43553\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43571\,
            I => \N__43550\
        );

    \I__9719\ : Span12Mux_v
    port map (
            O => \N__43566\,
            I => \N__43547\
        );

    \I__9718\ : Span4Mux_h
    port map (
            O => \N__43559\,
            I => \N__43542\
        );

    \I__9717\ : Span4Mux_h
    port map (
            O => \N__43556\,
            I => \N__43542\
        );

    \I__9716\ : Sp12to4
    port map (
            O => \N__43553\,
            I => \N__43539\
        );

    \I__9715\ : Span4Mux_h
    port map (
            O => \N__43550\,
            I => \N__43536\
        );

    \I__9714\ : Odrv12
    port map (
            O => \N__43547\,
            I => start_stop_c
        );

    \I__9713\ : Odrv4
    port map (
            O => \N__43542\,
            I => start_stop_c
        );

    \I__9712\ : Odrv12
    port map (
            O => \N__43539\,
            I => start_stop_c
        );

    \I__9711\ : Odrv4
    port map (
            O => \N__43536\,
            I => start_stop_c
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__43527\,
            I => \N__43524\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43521\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43518\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__43518\,
            I => \N__43515\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__43515\,
            I => \N__43509\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43506\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43503\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43512\,
            I => \N__43500\
        );

    \I__9702\ : Sp12to4
    port map (
            O => \N__43509\,
            I => \N__43495\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__43506\,
            I => \N__43495\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__43503\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__43500\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__9698\ : Odrv12
    port map (
            O => \N__43495\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__9697\ : CascadeMux
    port map (
            O => \N__43488\,
            I => \N__43485\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43482\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43482\,
            I => \N__43479\
        );

    \I__9694\ : Odrv4
    port map (
            O => \N__43479\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__9693\ : InMux
    port map (
            O => \N__43476\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__43473\,
            I => \N__43470\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43467\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43467\,
            I => \N__43463\
        );

    \I__9689\ : InMux
    port map (
            O => \N__43466\,
            I => \N__43458\
        );

    \I__9688\ : Sp12to4
    port map (
            O => \N__43463\,
            I => \N__43455\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43452\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43461\,
            I => \N__43449\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43458\,
            I => \N__43446\
        );

    \I__9684\ : Span12Mux_v
    port map (
            O => \N__43455\,
            I => \N__43443\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__43452\,
            I => \N__43440\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43449\,
            I => \N__43437\
        );

    \I__9681\ : Span4Mux_h
    port map (
            O => \N__43446\,
            I => \N__43434\
        );

    \I__9680\ : Odrv12
    port map (
            O => \N__43443\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__43440\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__9678\ : Odrv4
    port map (
            O => \N__43437\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__43434\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__9676\ : InMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__43422\,
            I => \N__43419\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__43419\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43416\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__9672\ : InMux
    port map (
            O => \N__43413\,
            I => \N__43410\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__43410\,
            I => \N__43407\
        );

    \I__9670\ : Span4Mux_v
    port map (
            O => \N__43407\,
            I => \N__43404\
        );

    \I__9669\ : Sp12to4
    port map (
            O => \N__43404\,
            I => \N__43399\
        );

    \I__9668\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43396\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43392\
        );

    \I__9666\ : Span12Mux_h
    port map (
            O => \N__43399\,
            I => \N__43389\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43386\
        );

    \I__9664\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43383\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__43392\,
            I => \N__43380\
        );

    \I__9662\ : Odrv12
    port map (
            O => \N__43389\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__9661\ : Odrv4
    port map (
            O => \N__43386\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__43383\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__9659\ : Odrv12
    port map (
            O => \N__43380\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43368\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43368\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43365\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__9655\ : CascadeMux
    port map (
            O => \N__43362\,
            I => \N__43359\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43355\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__43358\,
            I => \N__43352\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43355\,
            I => \N__43349\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43345\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__43349\,
            I => \N__43342\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__43348\,
            I => \N__43339\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43336\
        );

    \I__9647\ : Sp12to4
    port map (
            O => \N__43342\,
            I => \N__43332\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43329\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__43336\,
            I => \N__43326\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43323\
        );

    \I__9643\ : Span12Mux_h
    port map (
            O => \N__43332\,
            I => \N__43320\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__43329\,
            I => \N__43317\
        );

    \I__9641\ : Span4Mux_h
    port map (
            O => \N__43326\,
            I => \N__43314\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43323\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__9639\ : Odrv12
    port map (
            O => \N__43320\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__9638\ : Odrv4
    port map (
            O => \N__43317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__9637\ : Odrv4
    port map (
            O => \N__43314\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43302\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__43302\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43299\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__9633\ : CascadeMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__9632\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43290\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__9630\ : Span4Mux_h
    port map (
            O => \N__43287\,
            I => \N__43283\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43286\,
            I => \N__43279\
        );

    \I__9628\ : Span4Mux_v
    port map (
            O => \N__43283\,
            I => \N__43276\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43273\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43279\,
            I => \N__43269\
        );

    \I__9625\ : Span4Mux_h
    port map (
            O => \N__43276\,
            I => \N__43264\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__43273\,
            I => \N__43264\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43272\,
            I => \N__43261\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__43269\,
            I => \N__43256\
        );

    \I__9621\ : Span4Mux_h
    port map (
            O => \N__43264\,
            I => \N__43256\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__43261\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__43256\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__9618\ : InMux
    port map (
            O => \N__43251\,
            I => \N__43248\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__43248\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43245\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__9614\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43236\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43236\,
            I => \N__43233\
        );

    \I__9612\ : Span4Mux_v
    port map (
            O => \N__43233\,
            I => \N__43228\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__43232\,
            I => \N__43225\
        );

    \I__9610\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43222\
        );

    \I__9609\ : Span4Mux_h
    port map (
            O => \N__43228\,
            I => \N__43219\
        );

    \I__9608\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43215\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__43222\,
            I => \N__43212\
        );

    \I__9606\ : Span4Mux_h
    port map (
            O => \N__43219\,
            I => \N__43209\
        );

    \I__9605\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43206\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43203\
        );

    \I__9603\ : Span4Mux_v
    port map (
            O => \N__43212\,
            I => \N__43200\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__43209\,
            I => \N__43197\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43206\,
            I => \N__43190\
        );

    \I__9600\ : Span4Mux_v
    port map (
            O => \N__43203\,
            I => \N__43190\
        );

    \I__9599\ : Span4Mux_h
    port map (
            O => \N__43200\,
            I => \N__43190\
        );

    \I__9598\ : Odrv4
    port map (
            O => \N__43197\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9597\ : Odrv4
    port map (
            O => \N__43190\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__9596\ : CascadeMux
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__9595\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43179\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__43179\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43176\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__9592\ : CascadeMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__9591\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43162\
        );

    \I__9589\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43159\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43156\
        );

    \I__9587\ : Sp12to4
    port map (
            O => \N__43162\,
            I => \N__43152\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__43159\,
            I => \N__43147\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43156\,
            I => \N__43147\
        );

    \I__9584\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43144\
        );

    \I__9583\ : Span12Mux_v
    port map (
            O => \N__43152\,
            I => \N__43141\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__43147\,
            I => \N__43138\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43144\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9580\ : Odrv12
    port map (
            O => \N__43141\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9579\ : Odrv4
    port map (
            O => \N__43138\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__43131\,
            I => \N__43128\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__43122\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__9574\ : InMux
    port map (
            O => \N__43119\,
            I => \bfn_17_23_0_\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__43116\,
            I => \N__43113\
        );

    \I__9572\ : InMux
    port map (
            O => \N__43113\,
            I => \N__43110\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__9570\ : Span4Mux_v
    port map (
            O => \N__43107\,
            I => \N__43103\
        );

    \I__9569\ : InMux
    port map (
            O => \N__43106\,
            I => \N__43100\
        );

    \I__9568\ : Span4Mux_h
    port map (
            O => \N__43103\,
            I => \N__43097\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__43100\,
            I => \N__43093\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__43097\,
            I => \N__43089\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43096\,
            I => \N__43086\
        );

    \I__9564\ : Span4Mux_v
    port map (
            O => \N__43093\,
            I => \N__43083\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43092\,
            I => \N__43080\
        );

    \I__9562\ : Span4Mux_h
    port map (
            O => \N__43089\,
            I => \N__43077\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43086\,
            I => \N__43074\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__43083\,
            I => \N__43071\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__43080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__43077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__43074\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__43071\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9555\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43059\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43059\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__9553\ : InMux
    port map (
            O => \N__43056\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__9552\ : CascadeMux
    port map (
            O => \N__43053\,
            I => \N__43050\
        );

    \I__9551\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43047\,
            I => \N__43044\
        );

    \I__9549\ : Span4Mux_h
    port map (
            O => \N__43044\,
            I => \N__43041\
        );

    \I__9548\ : Span4Mux_h
    port map (
            O => \N__43041\,
            I => \N__43038\
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__43038\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__9546\ : InMux
    port map (
            O => \N__43035\,
            I => \N__43032\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__43032\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__9544\ : InMux
    port map (
            O => \N__43029\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__9543\ : CascadeMux
    port map (
            O => \N__43026\,
            I => \N__43023\
        );

    \I__9542\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__9540\ : Span4Mux_h
    port map (
            O => \N__43017\,
            I => \N__43014\
        );

    \I__9539\ : Span4Mux_h
    port map (
            O => \N__43014\,
            I => \N__43011\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__43011\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__9537\ : InMux
    port map (
            O => \N__43008\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__43005\,
            I => \N__43002\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__42999\,
            I => \N__42996\
        );

    \I__9533\ : Span4Mux_v
    port map (
            O => \N__42996\,
            I => \N__42993\
        );

    \I__9532\ : Sp12to4
    port map (
            O => \N__42993\,
            I => \N__42990\
        );

    \I__9531\ : Odrv12
    port map (
            O => \N__42990\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42987\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42984\,
            I => \N__42981\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__42981\,
            I => \N__42978\
        );

    \I__9527\ : Span4Mux_h
    port map (
            O => \N__42978\,
            I => \N__42974\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42971\
        );

    \I__9525\ : Span4Mux_v
    port map (
            O => \N__42974\,
            I => \N__42968\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42971\,
            I => \N__42965\
        );

    \I__9523\ : Span4Mux_h
    port map (
            O => \N__42968\,
            I => \N__42960\
        );

    \I__9522\ : Span4Mux_h
    port map (
            O => \N__42965\,
            I => \N__42960\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__42960\,
            I => \N__42955\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42952\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42949\
        );

    \I__9518\ : Odrv4
    port map (
            O => \N__42955\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__42949\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__42942\,
            I => \N__42939\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42936\,
            I => \N__42933\
        );

    \I__9512\ : Span4Mux_v
    port map (
            O => \N__42933\,
            I => \N__42930\
        );

    \I__9511\ : Span4Mux_h
    port map (
            O => \N__42930\,
            I => \N__42927\
        );

    \I__9510\ : Odrv4
    port map (
            O => \N__42927\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42924\,
            I => \N__42921\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42921\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42918\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__9506\ : CascadeMux
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__42906\,
            I => \N__42902\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42899\
        );

    \I__9501\ : Span4Mux_v
    port map (
            O => \N__42902\,
            I => \N__42894\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42899\,
            I => \N__42894\
        );

    \I__9499\ : Span4Mux_h
    port map (
            O => \N__42894\,
            I => \N__42889\
        );

    \I__9498\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42886\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42883\
        );

    \I__9496\ : Span4Mux_h
    port map (
            O => \N__42889\,
            I => \N__42880\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42886\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42883\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__42880\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__42873\,
            I => \N__42870\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42867\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42864\
        );

    \I__9489\ : Span4Mux_h
    port map (
            O => \N__42864\,
            I => \N__42861\
        );

    \I__9488\ : Span4Mux_h
    port map (
            O => \N__42861\,
            I => \N__42858\
        );

    \I__9487\ : Odrv4
    port map (
            O => \N__42858\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__9486\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42852\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42852\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42849\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__9483\ : CascadeMux
    port map (
            O => \N__42846\,
            I => \N__42843\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42840\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42837\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__42837\,
            I => \N__42832\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42836\,
            I => \N__42829\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42835\,
            I => \N__42826\
        );

    \I__9477\ : Sp12to4
    port map (
            O => \N__42832\,
            I => \N__42822\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42829\,
            I => \N__42819\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42826\,
            I => \N__42816\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42813\
        );

    \I__9473\ : Span12Mux_h
    port map (
            O => \N__42822\,
            I => \N__42810\
        );

    \I__9472\ : Span12Mux_h
    port map (
            O => \N__42819\,
            I => \N__42807\
        );

    \I__9471\ : Odrv4
    port map (
            O => \N__42816\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42813\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__9469\ : Odrv12
    port map (
            O => \N__42810\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__9468\ : Odrv12
    port map (
            O => \N__42807\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__42798\,
            I => \N__42795\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42792\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42792\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42789\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__9463\ : CascadeMux
    port map (
            O => \N__42786\,
            I => \N__42783\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42780\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42780\,
            I => \N__42777\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__42777\,
            I => \N__42773\
        );

    \I__9459\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42769\
        );

    \I__9458\ : Span4Mux_v
    port map (
            O => \N__42773\,
            I => \N__42766\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42763\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42769\,
            I => \N__42759\
        );

    \I__9455\ : Span4Mux_h
    port map (
            O => \N__42766\,
            I => \N__42754\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__42763\,
            I => \N__42754\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42751\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__42759\,
            I => \N__42746\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__42754\,
            I => \N__42746\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__42751\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__9449\ : Odrv4
    port map (
            O => \N__42746\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42738\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42738\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42735\,
            I => \bfn_17_22_0_\
        );

    \I__9445\ : CascadeMux
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42729\,
            I => \N__42726\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42726\,
            I => \N__42723\
        );

    \I__9442\ : Span4Mux_h
    port map (
            O => \N__42723\,
            I => \N__42720\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__42720\,
            I => \N__42714\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42719\,
            I => \N__42711\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42718\,
            I => \N__42708\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42705\
        );

    \I__9437\ : Span4Mux_h
    port map (
            O => \N__42714\,
            I => \N__42700\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42711\,
            I => \N__42700\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42708\,
            I => \N__42697\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42705\,
            I => \N__42694\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__42700\,
            I => \N__42691\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42697\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__42694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__42691\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__42684\,
            I => \N__42681\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__9426\ : Odrv4
    port map (
            O => \N__42675\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42672\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__9424\ : CascadeMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__9421\ : Span4Mux_v
    port map (
            O => \N__42660\,
            I => \N__42656\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42651\
        );

    \I__9419\ : Span4Mux_v
    port map (
            O => \N__42656\,
            I => \N__42648\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42645\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42642\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__42651\,
            I => \N__42639\
        );

    \I__9415\ : Span4Mux_h
    port map (
            O => \N__42648\,
            I => \N__42636\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42645\,
            I => \N__42633\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42642\,
            I => \N__42630\
        );

    \I__9412\ : Span4Mux_h
    port map (
            O => \N__42639\,
            I => \N__42623\
        );

    \I__9411\ : Span4Mux_h
    port map (
            O => \N__42636\,
            I => \N__42623\
        );

    \I__9410\ : Span4Mux_h
    port map (
            O => \N__42633\,
            I => \N__42623\
        );

    \I__9409\ : Odrv4
    port map (
            O => \N__42630\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__9408\ : Odrv4
    port map (
            O => \N__42623\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__9406\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42612\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__9404\ : Span4Mux_h
    port map (
            O => \N__42609\,
            I => \N__42606\
        );

    \I__9403\ : Span4Mux_h
    port map (
            O => \N__42606\,
            I => \N__42603\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__42603\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__9401\ : CascadeMux
    port map (
            O => \N__42600\,
            I => \N__42597\
        );

    \I__9400\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42594\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__42594\,
            I => \N__42591\
        );

    \I__9398\ : Span4Mux_v
    port map (
            O => \N__42591\,
            I => \N__42588\
        );

    \I__9397\ : Odrv4
    port map (
            O => \N__42588\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42585\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__42579\,
            I => \N__42576\
        );

    \I__9393\ : Span12Mux_v
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__9392\ : Odrv12
    port map (
            O => \N__42573\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__9391\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42565\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__42569\,
            I => \N__42562\
        );

    \I__9389\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42558\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42565\,
            I => \N__42555\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42562\,
            I => \N__42552\
        );

    \I__9386\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42549\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42558\,
            I => \N__42546\
        );

    \I__9384\ : Span4Mux_h
    port map (
            O => \N__42555\,
            I => \N__42543\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42538\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__42549\,
            I => \N__42538\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__42546\,
            I => \N__42535\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__42543\,
            I => \N__42532\
        );

    \I__9379\ : Span12Mux_h
    port map (
            O => \N__42538\,
            I => \N__42529\
        );

    \I__9378\ : Span4Mux_v
    port map (
            O => \N__42535\,
            I => \N__42524\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__42532\,
            I => \N__42524\
        );

    \I__9376\ : Odrv12
    port map (
            O => \N__42529\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__9375\ : Odrv4
    port map (
            O => \N__42524\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42516\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__42516\,
            I => \N__42513\
        );

    \I__9372\ : Span12Mux_s9_h
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__42510\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42507\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__9369\ : CascadeMux
    port map (
            O => \N__42504\,
            I => \N__42501\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42501\,
            I => \N__42498\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42498\,
            I => \N__42495\
        );

    \I__9366\ : Span4Mux_v
    port map (
            O => \N__42495\,
            I => \N__42492\
        );

    \I__9365\ : Span4Mux_h
    port map (
            O => \N__42492\,
            I => \N__42489\
        );

    \I__9364\ : Odrv4
    port map (
            O => \N__42489\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42486\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__9362\ : CascadeMux
    port map (
            O => \N__42483\,
            I => \N__42480\
        );

    \I__9361\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42477\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__42477\,
            I => \N__42474\
        );

    \I__9359\ : Span4Mux_h
    port map (
            O => \N__42474\,
            I => \N__42471\
        );

    \I__9358\ : Span4Mux_h
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__9357\ : Odrv4
    port map (
            O => \N__42468\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42465\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42453\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42450\
        );

    \I__9352\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42447\
        );

    \I__9351\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42444\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42441\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42450\,
            I => \N__42438\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42447\,
            I => \N__42433\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__42444\,
            I => \N__42433\
        );

    \I__9346\ : Span12Mux_h
    port map (
            O => \N__42441\,
            I => \N__42430\
        );

    \I__9345\ : Span4Mux_v
    port map (
            O => \N__42438\,
            I => \N__42425\
        );

    \I__9344\ : Span4Mux_v
    port map (
            O => \N__42433\,
            I => \N__42425\
        );

    \I__9343\ : Odrv12
    port map (
            O => \N__42430\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__42425\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__9341\ : CascadeMux
    port map (
            O => \N__42420\,
            I => \N__42417\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42414\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__42414\,
            I => \N__42411\
        );

    \I__9338\ : Span4Mux_h
    port map (
            O => \N__42411\,
            I => \N__42408\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__42405\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__9335\ : CascadeMux
    port map (
            O => \N__42402\,
            I => \N__42399\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42396\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42393\
        );

    \I__9332\ : Span4Mux_h
    port map (
            O => \N__42393\,
            I => \N__42390\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__42390\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42387\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__9329\ : CascadeMux
    port map (
            O => \N__42384\,
            I => \N__42381\
        );

    \I__9328\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__42378\,
            I => \N__42375\
        );

    \I__9326\ : Sp12to4
    port map (
            O => \N__42375\,
            I => \N__42370\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42366\
        );

    \I__9324\ : InMux
    port map (
            O => \N__42373\,
            I => \N__42363\
        );

    \I__9323\ : Span12Mux_h
    port map (
            O => \N__42370\,
            I => \N__42360\
        );

    \I__9322\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42357\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__42366\,
            I => \N__42354\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__42363\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9319\ : Odrv12
    port map (
            O => \N__42360\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__42357\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9317\ : Odrv4
    port map (
            O => \N__42354\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__9316\ : CascadeMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42342\,
            I => \N__42339\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__9312\ : Span4Mux_h
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__42330\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42324\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__42324\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42321\,
            I => \bfn_17_21_0_\
        );

    \I__9307\ : CascadeMux
    port map (
            O => \N__42318\,
            I => \N__42315\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42312\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42312\,
            I => \N__42309\
        );

    \I__9304\ : Span4Mux_h
    port map (
            O => \N__42309\,
            I => \N__42305\
        );

    \I__9303\ : InMux
    port map (
            O => \N__42308\,
            I => \N__42302\
        );

    \I__9302\ : Span4Mux_v
    port map (
            O => \N__42305\,
            I => \N__42296\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__42302\,
            I => \N__42296\
        );

    \I__9300\ : CascadeMux
    port map (
            O => \N__42301\,
            I => \N__42293\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__42296\,
            I => \N__42289\
        );

    \I__9298\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42286\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42292\,
            I => \N__42283\
        );

    \I__9296\ : Span4Mux_h
    port map (
            O => \N__42289\,
            I => \N__42280\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42286\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__42283\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__42280\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__42273\,
            I => \N__42270\
        );

    \I__9291\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42267\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__42267\,
            I => \N__42264\
        );

    \I__9289\ : Span4Mux_h
    port map (
            O => \N__42264\,
            I => \N__42261\
        );

    \I__9288\ : Span4Mux_h
    port map (
            O => \N__42261\,
            I => \N__42258\
        );

    \I__9287\ : Span4Mux_s0_h
    port map (
            O => \N__42258\,
            I => \N__42255\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42255\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__9285\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__42249\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42246\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__42243\,
            I => \N__42240\
        );

    \I__9281\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42237\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42237\,
            I => \N__42233\
        );

    \I__9279\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42230\
        );

    \I__9278\ : Span4Mux_v
    port map (
            O => \N__42233\,
            I => \N__42227\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__42230\,
            I => \N__42223\
        );

    \I__9276\ : Sp12to4
    port map (
            O => \N__42227\,
            I => \N__42219\
        );

    \I__9275\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42216\
        );

    \I__9274\ : Span12Mux_v
    port map (
            O => \N__42223\,
            I => \N__42213\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42210\
        );

    \I__9272\ : Span12Mux_h
    port map (
            O => \N__42219\,
            I => \N__42207\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__42216\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__9270\ : Odrv12
    port map (
            O => \N__42213\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__42210\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__9268\ : Odrv12
    port map (
            O => \N__42207\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__9267\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42195\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42195\,
            I => \N__42192\
        );

    \I__9265\ : Span4Mux_v
    port map (
            O => \N__42192\,
            I => \N__42188\
        );

    \I__9264\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42184\
        );

    \I__9263\ : Span4Mux_v
    port map (
            O => \N__42188\,
            I => \N__42181\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42187\,
            I => \N__42178\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__42184\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__42181\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__42178\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42165\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42165\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42165\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__9255\ : CascadeMux
    port map (
            O => \N__42162\,
            I => \N__42159\
        );

    \I__9254\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42156\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__42156\,
            I => \N__42153\
        );

    \I__9252\ : Span4Mux_h
    port map (
            O => \N__42153\,
            I => \N__42149\
        );

    \I__9251\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42146\
        );

    \I__9250\ : Sp12to4
    port map (
            O => \N__42149\,
            I => \N__42143\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__42146\,
            I => \N__42140\
        );

    \I__9248\ : Span12Mux_v
    port map (
            O => \N__42143\,
            I => \N__42137\
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__42140\,
            I => \phase_controller_inst2.stoper_hc.N_47\
        );

    \I__9246\ : Odrv12
    port map (
            O => \N__42137\,
            I => \phase_controller_inst2.stoper_hc.N_47\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42129\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__42129\,
            I => \N__42125\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42122\
        );

    \I__9242\ : Span4Mux_v
    port map (
            O => \N__42125\,
            I => \N__42119\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42122\,
            I => \N__42116\
        );

    \I__9240\ : Sp12to4
    port map (
            O => \N__42119\,
            I => \N__42112\
        );

    \I__9239\ : Span12Mux_v
    port map (
            O => \N__42116\,
            I => \N__42109\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42106\
        );

    \I__9237\ : Span12Mux_h
    port map (
            O => \N__42112\,
            I => \N__42103\
        );

    \I__9236\ : Span12Mux_v
    port map (
            O => \N__42109\,
            I => \N__42098\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42098\
        );

    \I__9234\ : Span12Mux_v
    port map (
            O => \N__42103\,
            I => \N__42093\
        );

    \I__9233\ : Span12Mux_h
    port map (
            O => \N__42098\,
            I => \N__42093\
        );

    \I__9232\ : Odrv12
    port map (
            O => \N__42093\,
            I => il_max_comp2_c
        );

    \I__9231\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42084\
        );

    \I__9230\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42084\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__42084\,
            I => \N__42080\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42077\
        );

    \I__9227\ : Span4Mux_v
    port map (
            O => \N__42080\,
            I => \N__42074\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42077\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__42074\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42069\,
            I => \N__42065\
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__42068\,
            I => \N__42061\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42065\,
            I => \N__42058\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42053\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42061\,
            I => \N__42053\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__42058\,
            I => \N__42050\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__42053\,
            I => \N__42046\
        );

    \I__9217\ : Span4Mux_v
    port map (
            O => \N__42050\,
            I => \N__42042\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42039\
        );

    \I__9215\ : Span4Mux_v
    port map (
            O => \N__42046\,
            I => \N__42036\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42033\
        );

    \I__9213\ : Span4Mux_v
    port map (
            O => \N__42042\,
            I => \N__42030\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__42025\
        );

    \I__9211\ : Span4Mux_h
    port map (
            O => \N__42036\,
            I => \N__42025\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__42033\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__42030\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__42025\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__9207\ : InMux
    port map (
            O => \N__42018\,
            I => \N__42014\
        );

    \I__9206\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42011\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__42014\,
            I => \N__42006\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__42011\,
            I => \N__42006\
        );

    \I__9203\ : Span4Mux_v
    port map (
            O => \N__42006\,
            I => \N__42000\
        );

    \I__9202\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41993\
        );

    \I__9201\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41993\
        );

    \I__9200\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41993\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__42000\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41993\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41985\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41985\,
            I => \N__41981\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41978\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__41981\,
            I => \N__41975\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__41978\,
            I => \N__41972\
        );

    \I__9192\ : Span4Mux_v
    port map (
            O => \N__41975\,
            I => \N__41969\
        );

    \I__9191\ : Span4Mux_h
    port map (
            O => \N__41972\,
            I => \N__41964\
        );

    \I__9190\ : Span4Mux_v
    port map (
            O => \N__41969\,
            I => \N__41964\
        );

    \I__9189\ : Odrv4
    port map (
            O => \N__41964\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__41949\,
            I => \phase_controller_inst2.stoper_hc.mZ0Z16\
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__41946\,
            I => \N__41943\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__9180\ : Span4Mux_h
    port map (
            O => \N__41937\,
            I => \N__41934\
        );

    \I__9179\ : Sp12to4
    port map (
            O => \N__41934\,
            I => \N__41931\
        );

    \I__9178\ : Span12Mux_v
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__9177\ : Odrv12
    port map (
            O => \N__41928\,
            I => \phase_controller_inst2.stoper_hc.m28_ns_1\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41925\,
            I => \N__41919\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41924\,
            I => \N__41919\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41919\,
            I => \N__41915\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41918\,
            I => \N__41912\
        );

    \I__9172\ : Span4Mux_h
    port map (
            O => \N__41915\,
            I => \N__41909\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41912\,
            I => \N__41905\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__41909\,
            I => \N__41902\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41908\,
            I => \N__41899\
        );

    \I__9168\ : Span12Mux_h
    port map (
            O => \N__41905\,
            I => \N__41896\
        );

    \I__9167\ : Span4Mux_v
    port map (
            O => \N__41902\,
            I => \N__41893\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41899\,
            I => \N__41888\
        );

    \I__9165\ : Span12Mux_v
    port map (
            O => \N__41896\,
            I => \N__41885\
        );

    \I__9164\ : Span4Mux_v
    port map (
            O => \N__41893\,
            I => \N__41882\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41879\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41876\
        );

    \I__9161\ : Span4Mux_h
    port map (
            O => \N__41888\,
            I => \N__41873\
        );

    \I__9160\ : Odrv12
    port map (
            O => \N__41885\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__41882\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41879\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41876\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__41873\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41859\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41859\,
            I => \N__41853\
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__41858\,
            I => \N__41850\
        );

    \I__9152\ : CascadeMux
    port map (
            O => \N__41857\,
            I => \N__41847\
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__41856\,
            I => \N__41844\
        );

    \I__9150\ : Span4Mux_h
    port map (
            O => \N__41853\,
            I => \N__41840\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41837\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41832\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41844\,
            I => \N__41832\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41829\
        );

    \I__9145\ : Sp12to4
    port map (
            O => \N__41840\,
            I => \N__41820\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__41837\,
            I => \N__41820\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41832\,
            I => \N__41820\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__41829\,
            I => \N__41820\
        );

    \I__9141\ : Span12Mux_s6_v
    port map (
            O => \N__41820\,
            I => \N__41816\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41819\,
            I => \N__41813\
        );

    \I__9139\ : Span12Mux_v
    port map (
            O => \N__41816\,
            I => \N__41810\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41813\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9137\ : Odrv12
    port map (
            O => \N__41810\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9136\ : CascadeMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41799\,
            I => \N__41796\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__41796\,
            I => \N__41791\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41795\,
            I => \N__41787\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__41794\,
            I => \N__41784\
        );

    \I__9130\ : Span4Mux_v
    port map (
            O => \N__41791\,
            I => \N__41781\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41778\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41787\,
            I => \N__41774\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41771\
        );

    \I__9126\ : Span4Mux_h
    port map (
            O => \N__41781\,
            I => \N__41768\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41778\,
            I => \N__41765\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41762\
        );

    \I__9123\ : Span12Mux_h
    port map (
            O => \N__41774\,
            I => \N__41759\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41771\,
            I => \N__41756\
        );

    \I__9121\ : Span4Mux_h
    port map (
            O => \N__41768\,
            I => \N__41751\
        );

    \I__9120\ : Span4Mux_v
    port map (
            O => \N__41765\,
            I => \N__41751\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__41762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__9118\ : Odrv12
    port map (
            O => \N__41759\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__9117\ : Odrv4
    port map (
            O => \N__41756\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__9116\ : Odrv4
    port map (
            O => \N__41751\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__9115\ : CascadeMux
    port map (
            O => \N__41742\,
            I => \N__41739\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41735\
        );

    \I__9113\ : CascadeMux
    port map (
            O => \N__41738\,
            I => \N__41732\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__41735\,
            I => \N__41729\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41732\,
            I => \N__41726\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__41729\,
            I => \N__41723\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41726\,
            I => \N__41720\
        );

    \I__9108\ : Span4Mux_h
    port map (
            O => \N__41723\,
            I => \N__41717\
        );

    \I__9107\ : Span4Mux_h
    port map (
            O => \N__41720\,
            I => \N__41714\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__41717\,
            I => \N__41711\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__41714\,
            I => \N__41708\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__41711\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__41708\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__9102\ : CascadeMux
    port map (
            O => \N__41703\,
            I => \N__41700\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41694\
        );

    \I__9099\ : Span4Mux_v
    port map (
            O => \N__41694\,
            I => \N__41689\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41686\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41683\
        );

    \I__9096\ : Sp12to4
    port map (
            O => \N__41689\,
            I => \N__41680\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41686\,
            I => \N__41677\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41683\,
            I => \N__41672\
        );

    \I__9093\ : Span12Mux_h
    port map (
            O => \N__41680\,
            I => \N__41672\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__41677\,
            I => \N__41669\
        );

    \I__9091\ : Odrv12
    port map (
            O => \N__41672\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__9090\ : Odrv4
    port map (
            O => \N__41669\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__9089\ : CascadeMux
    port map (
            O => \N__41664\,
            I => \N__41661\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41658\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41655\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__41655\,
            I => \N__41652\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__41652\,
            I => \N__41649\
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__41649\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41640\
        );

    \I__9081\ : Span4Mux_v
    port map (
            O => \N__41640\,
            I => \N__41637\
        );

    \I__9080\ : Odrv4
    port map (
            O => \N__41637\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41634\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__9078\ : CascadeMux
    port map (
            O => \N__41631\,
            I => \N__41628\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41628\,
            I => \N__41624\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41627\,
            I => \N__41621\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41624\,
            I => \N__41618\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41621\,
            I => \N__41615\
        );

    \I__9073\ : Span4Mux_h
    port map (
            O => \N__41618\,
            I => \N__41610\
        );

    \I__9072\ : Span4Mux_h
    port map (
            O => \N__41615\,
            I => \N__41607\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41604\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41601\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__41610\,
            I => \N__41596\
        );

    \I__9068\ : Span4Mux_h
    port map (
            O => \N__41607\,
            I => \N__41596\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__41604\,
            I => \N__41591\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__41601\,
            I => \N__41591\
        );

    \I__9065\ : Odrv4
    port map (
            O => \N__41596\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__9064\ : Odrv12
    port map (
            O => \N__41591\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__41586\,
            I => \N__41583\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41580\,
            I => \N__41577\
        );

    \I__9060\ : Span4Mux_h
    port map (
            O => \N__41577\,
            I => \N__41574\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__41574\,
            I => \N__41571\
        );

    \I__9058\ : Odrv4
    port map (
            O => \N__41571\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41565\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__41565\,
            I => \N__41562\
        );

    \I__9055\ : Span12Mux_s11_h
    port map (
            O => \N__41562\,
            I => \N__41559\
        );

    \I__9054\ : Odrv12
    port map (
            O => \N__41559\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41556\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__9052\ : CascadeMux
    port map (
            O => \N__41553\,
            I => \N__41549\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41544\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41544\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__41544\,
            I => \N__41541\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__41541\,
            I => \N__41537\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41540\,
            I => \N__41534\
        );

    \I__9046\ : Span4Mux_h
    port map (
            O => \N__41537\,
            I => \N__41531\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__41534\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__9044\ : Odrv4
    port map (
            O => \N__41531\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41526\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41523\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41520\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__41517\,
            I => \N__41512\
        );

    \I__9039\ : InMux
    port map (
            O => \N__41516\,
            I => \N__41509\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41504\
        );

    \I__9037\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41504\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__41509\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__41504\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__9034\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41494\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41489\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41489\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41494\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41489\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41480\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41477\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41480\,
            I => \N__41473\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41477\,
            I => \N__41470\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41467\
        );

    \I__9024\ : Span4Mux_v
    port map (
            O => \N__41473\,
            I => \N__41464\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__41470\,
            I => \N__41461\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41467\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__41464\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9020\ : Odrv4
    port map (
            O => \N__41461\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9019\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41448\
        );

    \I__9018\ : InMux
    port map (
            O => \N__41453\,
            I => \N__41448\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__41448\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__9016\ : CascadeMux
    port map (
            O => \N__41445\,
            I => \N__41441\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41437\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41441\,
            I => \N__41432\
        );

    \I__9013\ : InMux
    port map (
            O => \N__41440\,
            I => \N__41432\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__41437\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41432\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__9010\ : CascadeMux
    port map (
            O => \N__41427\,
            I => \N__41424\
        );

    \I__9009\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41418\
        );

    \I__9008\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41418\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__41418\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41410\
        );

    \I__9005\ : InMux
    port map (
            O => \N__41414\,
            I => \N__41405\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41405\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__41410\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__41405\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__9001\ : CascadeMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__9000\ : InMux
    port map (
            O => \N__41397\,
            I => \N__41391\
        );

    \I__8999\ : InMux
    port map (
            O => \N__41396\,
            I => \N__41391\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41391\,
            I => \N__41387\
        );

    \I__8997\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41384\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__41387\,
            I => \N__41381\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41384\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__41381\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8993\ : InMux
    port map (
            O => \N__41376\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41366\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41366\
        );

    \I__8990\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41363\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41360\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41363\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8987\ : Odrv4
    port map (
            O => \N__41360\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41355\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41352\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__8984\ : InMux
    port map (
            O => \N__41349\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41339\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41339\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41336\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__41339\,
            I => \N__41333\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41336\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__41333\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41328\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41320\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41315\
        );

    \I__8974\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41315\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__41320\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__41315\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41310\,
            I => \bfn_17_17_0_\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41307\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41304\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41295\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41300\,
            I => \N__41295\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__41295\,
            I => \N__41292\
        );

    \I__8965\ : Span4Mux_v
    port map (
            O => \N__41292\,
            I => \N__41288\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41291\,
            I => \N__41285\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__41288\,
            I => \N__41282\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__41285\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__41282\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8960\ : InMux
    port map (
            O => \N__41277\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41274\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41271\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41268\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41265\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41262\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41259\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41256\,
            I => \bfn_17_16_0_\
        );

    \I__8952\ : InMux
    port map (
            O => \N__41253\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41250\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41247\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__41244\,
            I => \N__41240\
        );

    \I__8948\ : CascadeMux
    port map (
            O => \N__41243\,
            I => \N__41237\
        );

    \I__8947\ : InMux
    port map (
            O => \N__41240\,
            I => \N__41232\
        );

    \I__8946\ : InMux
    port map (
            O => \N__41237\,
            I => \N__41232\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__41232\,
            I => \phase_controller_inst2.stoper_hc.N_265_i\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41229\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41226\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41223\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__8941\ : InMux
    port map (
            O => \N__41220\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41217\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41214\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__8938\ : InMux
    port map (
            O => \N__41211\,
            I => \bfn_17_15_0_\
        );

    \I__8937\ : InMux
    port map (
            O => \N__41208\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__8936\ : InMux
    port map (
            O => \N__41205\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41202\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__8934\ : InMux
    port map (
            O => \N__41199\,
            I => \bfn_17_13_0_\
        );

    \I__8933\ : InMux
    port map (
            O => \N__41196\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__8932\ : InMux
    port map (
            O => \N__41193\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41190\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__8930\ : InMux
    port map (
            O => \N__41187\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__8929\ : InMux
    port map (
            O => \N__41184\,
            I => \N__41168\
        );

    \I__8928\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41168\
        );

    \I__8927\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41168\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41168\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41143\
        );

    \I__8924\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41143\
        );

    \I__8923\ : InMux
    port map (
            O => \N__41178\,
            I => \N__41143\
        );

    \I__8922\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41143\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__41168\,
            I => \N__41134\
        );

    \I__8920\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41125\
        );

    \I__8919\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41125\
        );

    \I__8918\ : InMux
    port map (
            O => \N__41165\,
            I => \N__41125\
        );

    \I__8917\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41125\
        );

    \I__8916\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41116\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41116\
        );

    \I__8914\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41116\
        );

    \I__8913\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41116\
        );

    \I__8912\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41107\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41107\
        );

    \I__8910\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41107\
        );

    \I__8909\ : InMux
    port map (
            O => \N__41156\,
            I => \N__41107\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41155\,
            I => \N__41098\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41098\
        );

    \I__8906\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41098\
        );

    \I__8905\ : InMux
    port map (
            O => \N__41152\,
            I => \N__41098\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41095\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41090\
        );

    \I__8902\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41090\
        );

    \I__8901\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41081\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41081\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41081\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41081\
        );

    \I__8897\ : Span4Mux_v
    port map (
            O => \N__41134\,
            I => \N__41078\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__41125\,
            I => \N__41069\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41116\,
            I => \N__41069\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41107\,
            I => \N__41069\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41098\,
            I => \N__41069\
        );

    \I__8892\ : Span4Mux_h
    port map (
            O => \N__41095\,
            I => \N__41066\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41090\,
            I => \N__41057\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41081\,
            I => \N__41057\
        );

    \I__8889\ : Span4Mux_h
    port map (
            O => \N__41078\,
            I => \N__41057\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__41069\,
            I => \N__41057\
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__41066\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8886\ : Odrv4
    port map (
            O => \N__41057\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8885\ : InMux
    port map (
            O => \N__41052\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__8884\ : CEMux
    port map (
            O => \N__41049\,
            I => \N__41045\
        );

    \I__8883\ : CEMux
    port map (
            O => \N__41048\,
            I => \N__41042\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__41045\,
            I => \N__41037\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41034\
        );

    \I__8880\ : CEMux
    port map (
            O => \N__41041\,
            I => \N__41031\
        );

    \I__8879\ : CEMux
    port map (
            O => \N__41040\,
            I => \N__41028\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__41037\,
            I => \N__41025\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__41034\,
            I => \N__41022\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__41031\,
            I => \N__41019\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41016\
        );

    \I__8874\ : Span4Mux_v
    port map (
            O => \N__41025\,
            I => \N__41013\
        );

    \I__8873\ : Span4Mux_v
    port map (
            O => \N__41022\,
            I => \N__41010\
        );

    \I__8872\ : Span4Mux_h
    port map (
            O => \N__41019\,
            I => \N__41007\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__41016\,
            I => \N__41004\
        );

    \I__8870\ : Odrv4
    port map (
            O => \N__41013\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__41010\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__41007\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__8867\ : Odrv4
    port map (
            O => \N__41004\,
            I => \delay_measurement_inst.delay_hc_timer.N_342_i\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40995\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40992\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40989\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40986\,
            I => \bfn_17_12_0_\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40983\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40980\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__8860\ : InMux
    port map (
            O => \N__40977\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40974\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__8858\ : InMux
    port map (
            O => \N__40971\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40968\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40965\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40962\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__8854\ : InMux
    port map (
            O => \N__40959\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__8853\ : InMux
    port map (
            O => \N__40956\,
            I => \bfn_17_11_0_\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40953\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40950\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40947\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40944\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__8848\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40935\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40940\,
            I => \N__40935\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__40935\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40932\,
            I => \N__40929\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40929\,
            I => \N__40925\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40921\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__40925\,
            I => \N__40918\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40924\,
            I => \N__40915\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40921\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__40918\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__40915\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__40908\,
            I => \N__40905\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40902\,
            I => \N__40899\
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__40899\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40890\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40890\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40890\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40881\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40881\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40877\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40874\
        );

    \I__8826\ : Span4Mux_h
    port map (
            O => \N__40877\,
            I => \N__40871\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__40874\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8824\ : Odrv4
    port map (
            O => \N__40871\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8823\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40860\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40860\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40860\,
            I => \N__40856\
        );

    \I__8820\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40853\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__40856\,
            I => \N__40850\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40853\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__40850\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40842\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__40839\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40836\,
            I => \bfn_17_10_0_\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40833\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40830\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40827\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40821\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40821\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40812\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40817\,
            I => \N__40812\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40812\,
            I => \N__40808\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40811\,
            I => \N__40805\
        );

    \I__8803\ : Span4Mux_v
    port map (
            O => \N__40808\,
            I => \N__40802\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40805\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__40802\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__8800\ : CascadeMux
    port map (
            O => \N__40797\,
            I => \N__40792\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__40796\,
            I => \N__40789\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40786\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40783\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40789\,
            I => \N__40780\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__40786\,
            I => \N__40773\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40773\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40780\,
            I => \N__40773\
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__40773\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40767\,
            I => \N__40764\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40764\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40761\,
            I => \N__40755\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40755\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40755\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40752\,
            I => \N__40749\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40749\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40743\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40740\
        );

    \I__8781\ : Span4Mux_v
    port map (
            O => \N__40740\,
            I => \N__40737\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__40737\,
            I => \N__40733\
        );

    \I__8779\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40730\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__40733\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40730\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__8776\ : CascadeMux
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40722\,
            I => \N__40719\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__40719\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__40713\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40707\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__40707\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__8769\ : CascadeMux
    port map (
            O => \N__40704\,
            I => \N__40701\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40698\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40698\,
            I => \N__40695\
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__40695\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__40692\,
            I => \N__40687\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40684\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40679\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40679\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40684\,
            I => \N__40674\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__40679\,
            I => \N__40674\
        );

    \I__8759\ : Odrv4
    port map (
            O => \N__40674\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__40671\,
            I => \N__40666\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40663\
        );

    \I__8756\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40658\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40658\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40663\,
            I => \N__40653\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40653\
        );

    \I__8752\ : Odrv4
    port map (
            O => \N__40653\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40647\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40647\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40644\,
            I => \N__40639\
        );

    \I__8748\ : CascadeMux
    port map (
            O => \N__40643\,
            I => \N__40636\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40642\,
            I => \N__40632\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40628\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40625\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40622\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40632\,
            I => \N__40619\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40616\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__40628\,
            I => \N__40610\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40625\,
            I => \N__40610\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40622\,
            I => \N__40603\
        );

    \I__8738\ : Span4Mux_s2_v
    port map (
            O => \N__40619\,
            I => \N__40603\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__40616\,
            I => \N__40603\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40600\
        );

    \I__8735\ : Span4Mux_h
    port map (
            O => \N__40610\,
            I => \N__40597\
        );

    \I__8734\ : Span4Mux_h
    port map (
            O => \N__40603\,
            I => \N__40594\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40600\,
            I => \phase_controller_inst1.stoper_hc.hc_time_passed\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__40597\,
            I => \phase_controller_inst1.stoper_hc.hc_time_passed\
        );

    \I__8731\ : Odrv4
    port map (
            O => \N__40594\,
            I => \phase_controller_inst1.stoper_hc.hc_time_passed\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40583\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40580\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40583\,
            I => \phase_controller_inst1.stoper_hc.N_45\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40580\,
            I => \phase_controller_inst1.stoper_hc.N_45\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40571\
        );

    \I__8725\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40567\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40571\,
            I => \N__40564\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40561\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__40567\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8721\ : Odrv4
    port map (
            O => \N__40564\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__40561\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8719\ : CascadeMux
    port map (
            O => \N__40554\,
            I => \N__40547\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40553\,
            I => \N__40544\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40539\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40539\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40536\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40533\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40544\,
            I => \N__40530\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40539\,
            I => \N__40527\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40536\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__40533\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__40530\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__40527\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40513\
        );

    \I__8706\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40508\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40516\,
            I => \N__40505\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__40513\,
            I => \N__40502\
        );

    \I__8703\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40497\
        );

    \I__8702\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40497\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__40508\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__40505\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__40502\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40497\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__8697\ : CascadeMux
    port map (
            O => \N__40488\,
            I => \N__40483\
        );

    \I__8696\ : CascadeMux
    port map (
            O => \N__40487\,
            I => \N__40480\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40477\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40474\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40471\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__40477\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40474\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40471\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40460\
        );

    \I__8688\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40457\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__40460\,
            I => \N__40454\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40457\,
            I => \N__40451\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__40454\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8684\ : Odrv12
    port map (
            O => \N__40451\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40443\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40443\,
            I => \phase_controller_inst1.stoper_hc.N_46\
        );

    \I__8681\ : CascadeMux
    port map (
            O => \N__40440\,
            I => \phase_controller_inst1.stoper_hc.N_46_cascade_\
        );

    \I__8680\ : CEMux
    port map (
            O => \N__40437\,
            I => \N__40434\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40431\
        );

    \I__8678\ : Odrv4
    port map (
            O => \N__40431\,
            I => \phase_controller_inst1.stoper_hc.N_46_0\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__40428\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__8676\ : CascadeMux
    port map (
            O => \N__40425\,
            I => \current_shift_inst.PI_CTRL.N_287_cascade_\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40419\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__40419\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__8673\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40413\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__40413\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__40410\,
            I => \N__40407\
        );

    \I__8670\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40402\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40399\
        );

    \I__8668\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40396\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__40402\,
            I => \N__40391\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40399\,
            I => \N__40391\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__40396\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__40391\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8663\ : InMux
    port map (
            O => \N__40386\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40383\,
            I => \N__40376\
        );

    \I__8661\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40376\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40381\,
            I => \N__40373\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__40376\,
            I => \N__40370\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__40373\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8657\ : Odrv4
    port map (
            O => \N__40370\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8656\ : InMux
    port map (
            O => \N__40365\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40358\
        );

    \I__8654\ : InMux
    port map (
            O => \N__40361\,
            I => \N__40355\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__40358\,
            I => \N__40352\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__40355\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__40352\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8650\ : InMux
    port map (
            O => \N__40347\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40344\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40338\,
            I => \N__40334\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40337\,
            I => \N__40331\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__40334\,
            I => \N__40328\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40331\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__40328\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8642\ : CEMux
    port map (
            O => \N__40323\,
            I => \N__40319\
        );

    \I__8641\ : CEMux
    port map (
            O => \N__40322\,
            I => \N__40316\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__40319\,
            I => \N__40311\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40316\,
            I => \N__40308\
        );

    \I__8638\ : CEMux
    port map (
            O => \N__40315\,
            I => \N__40305\
        );

    \I__8637\ : CEMux
    port map (
            O => \N__40314\,
            I => \N__40302\
        );

    \I__8636\ : Span4Mux_v
    port map (
            O => \N__40311\,
            I => \N__40299\
        );

    \I__8635\ : Span4Mux_h
    port map (
            O => \N__40308\,
            I => \N__40296\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__40305\,
            I => \N__40291\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40302\,
            I => \N__40291\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__40299\,
            I => \current_shift_inst.timer_s1.N_340_i\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__40296\,
            I => \current_shift_inst.timer_s1.N_340_i\
        );

    \I__8630\ : Odrv4
    port map (
            O => \N__40291\,
            I => \current_shift_inst.timer_s1.N_340_i\
        );

    \I__8629\ : CascadeMux
    port map (
            O => \N__40284\,
            I => \N__40281\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40281\,
            I => \N__40275\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40275\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__40275\,
            I => \N__40272\
        );

    \I__8625\ : Span4Mux_v
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__40269\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__40266\,
            I => \N__40262\
        );

    \I__8622\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40257\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40257\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__8619\ : Odrv12
    port map (
            O => \N__40254\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__40251\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40245\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__40245\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40242\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__8614\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40232\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40232\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40229\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40226\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40229\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__40226\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40221\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40211\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40211\
        );

    \I__8605\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40208\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__40211\,
            I => \N__40205\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40208\,
            I => \N__40200\
        );

    \I__8602\ : Span4Mux_h
    port map (
            O => \N__40205\,
            I => \N__40200\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40200\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__8600\ : InMux
    port map (
            O => \N__40197\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__40194\,
            I => \N__40190\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40186\
        );

    \I__8597\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40183\
        );

    \I__8596\ : InMux
    port map (
            O => \N__40189\,
            I => \N__40180\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40186\,
            I => \N__40175\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40183\,
            I => \N__40175\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__40180\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__40175\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40170\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__8590\ : CascadeMux
    port map (
            O => \N__40167\,
            I => \N__40163\
        );

    \I__8589\ : InMux
    port map (
            O => \N__40166\,
            I => \N__40159\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40156\
        );

    \I__8587\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40153\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__40159\,
            I => \N__40148\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40156\,
            I => \N__40148\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__40153\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__40148\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40143\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__8581\ : CascadeMux
    port map (
            O => \N__40140\,
            I => \N__40136\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__40139\,
            I => \N__40133\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40136\,
            I => \N__40127\
        );

    \I__8578\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40127\
        );

    \I__8577\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40124\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__40127\,
            I => \N__40121\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40124\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__40121\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40116\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__40113\,
            I => \N__40109\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__40112\,
            I => \N__40106\
        );

    \I__8570\ : InMux
    port map (
            O => \N__40109\,
            I => \N__40100\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40106\,
            I => \N__40100\
        );

    \I__8568\ : InMux
    port map (
            O => \N__40105\,
            I => \N__40097\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__40097\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__40094\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8564\ : InMux
    port map (
            O => \N__40089\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__40086\,
            I => \N__40083\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40078\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40075\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40072\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__40078\,
            I => \N__40067\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40075\,
            I => \N__40067\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__40072\,
            I => \N__40062\
        );

    \I__8556\ : Span4Mux_v
    port map (
            O => \N__40067\,
            I => \N__40062\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__40062\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40059\,
            I => \bfn_16_17_0_\
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__40056\,
            I => \N__40053\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40053\,
            I => \N__40049\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40046\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40049\,
            I => \N__40040\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__40046\,
            I => \N__40040\
        );

    \I__8548\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40037\
        );

    \I__8547\ : Span4Mux_v
    port map (
            O => \N__40040\,
            I => \N__40034\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__40037\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__40034\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8544\ : InMux
    port map (
            O => \N__40029\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__40026\,
            I => \N__40022\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__40025\,
            I => \N__40019\
        );

    \I__8541\ : InMux
    port map (
            O => \N__40022\,
            I => \N__40016\
        );

    \I__8540\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40012\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__40016\,
            I => \N__40009\
        );

    \I__8538\ : InMux
    port map (
            O => \N__40015\,
            I => \N__40006\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__40012\,
            I => \N__40003\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__40009\,
            I => \N__40000\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__40006\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8534\ : Odrv12
    port map (
            O => \N__40003\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__40000\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39993\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39983\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39983\
        );

    \I__8529\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39980\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__39983\,
            I => \N__39977\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__39980\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__39977\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39972\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39969\,
            I => \N__39962\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39968\,
            I => \N__39962\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39967\,
            I => \N__39959\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39962\,
            I => \N__39956\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__39959\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8519\ : Odrv12
    port map (
            O => \N__39956\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39951\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__39948\,
            I => \N__39944\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39947\,
            I => \N__39940\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39937\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39943\,
            I => \N__39934\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39940\,
            I => \N__39929\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39937\,
            I => \N__39929\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__39934\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8510\ : Odrv4
    port map (
            O => \N__39929\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39924\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__39921\,
            I => \N__39917\
        );

    \I__8507\ : CascadeMux
    port map (
            O => \N__39920\,
            I => \N__39914\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39908\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39908\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39905\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39908\,
            I => \N__39902\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__39905\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8501\ : Odrv4
    port map (
            O => \N__39902\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8500\ : InMux
    port map (
            O => \N__39897\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__8499\ : CascadeMux
    port map (
            O => \N__39894\,
            I => \N__39890\
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__39893\,
            I => \N__39887\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39881\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39881\
        );

    \I__8495\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39878\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__39881\,
            I => \N__39875\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__39878\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8492\ : Odrv4
    port map (
            O => \N__39875\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39870\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39867\,
            I => \N__39860\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39866\,
            I => \N__39860\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39865\,
            I => \N__39857\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39860\,
            I => \N__39854\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39857\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__39854\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39849\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__8483\ : CascadeMux
    port map (
            O => \N__39846\,
            I => \N__39843\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39843\,
            I => \N__39838\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39835\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39832\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39827\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__39835\,
            I => \N__39827\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39832\,
            I => \N__39822\
        );

    \I__8476\ : Span4Mux_v
    port map (
            O => \N__39827\,
            I => \N__39822\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__39822\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39819\,
            I => \bfn_16_16_0_\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__39816\,
            I => \N__39812\
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__39815\,
            I => \N__39809\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39806\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39803\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39806\,
            I => \N__39799\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39796\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39793\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__39799\,
            I => \N__39788\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__39796\,
            I => \N__39788\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__39793\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__39788\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39783\,
            I => \N__39779\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__39782\,
            I => \N__39776\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39779\,
            I => \N__39773\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39769\
        );

    \I__8458\ : Span4Mux_h
    port map (
            O => \N__39773\,
            I => \N__39766\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39763\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__39769\,
            I => \N__39760\
        );

    \I__8455\ : Odrv4
    port map (
            O => \N__39766\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39763\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8453\ : Odrv12
    port map (
            O => \N__39760\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39753\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39743\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39749\,
            I => \N__39743\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39740\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39743\,
            I => \N__39737\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39740\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8446\ : Odrv12
    port map (
            O => \N__39737\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39732\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39722\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39722\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39727\,
            I => \N__39719\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39722\,
            I => \N__39716\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39719\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8439\ : Odrv12
    port map (
            O => \N__39716\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39711\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__39708\,
            I => \N__39704\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__39707\,
            I => \N__39701\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39695\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39701\,
            I => \N__39695\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39700\,
            I => \N__39692\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39695\,
            I => \N__39689\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39692\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8430\ : Odrv4
    port map (
            O => \N__39689\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39684\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__39681\,
            I => \N__39677\
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__39680\,
            I => \N__39674\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39668\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39668\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39665\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__39668\,
            I => \N__39662\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39665\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8421\ : Odrv4
    port map (
            O => \N__39662\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39657\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39647\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39647\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39644\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39647\,
            I => \N__39641\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39644\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__39641\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39636\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39626\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39626\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39623\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__39626\,
            I => \N__39620\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__39623\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__39620\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8406\ : InMux
    port map (
            O => \N__39615\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__39612\,
            I => \N__39608\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__39611\,
            I => \N__39605\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39601\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39598\
        );

    \I__8401\ : InMux
    port map (
            O => \N__39604\,
            I => \N__39595\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__39601\,
            I => \N__39590\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39598\,
            I => \N__39590\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__39595\,
            I => \N__39585\
        );

    \I__8397\ : Span4Mux_v
    port map (
            O => \N__39590\,
            I => \N__39585\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__39585\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39582\,
            I => \bfn_16_15_0_\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39574\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39578\,
            I => \N__39571\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39568\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__39574\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__39571\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__39568\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39556\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39560\,
            I => \N__39553\
        );

    \I__8386\ : InMux
    port map (
            O => \N__39559\,
            I => \N__39550\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__39556\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39553\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__39550\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__8382\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__39540\,
            I => \N__39536\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39532\
        );

    \I__8379\ : Span4Mux_h
    port map (
            O => \N__39536\,
            I => \N__39529\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39526\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__39532\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8376\ : Odrv4
    port map (
            O => \N__39529\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39526\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39514\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39511\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39508\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39514\,
            I => \N__39505\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__39511\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39508\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8368\ : Odrv4
    port map (
            O => \N__39505\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39492\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39492\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__39492\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__39489\,
            I => \N__39486\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39480\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39480\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__39480\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39473\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39469\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39473\,
            I => \N__39466\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39463\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39469\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__8355\ : Odrv4
    port map (
            O => \N__39466\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__39463\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39452\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__39455\,
            I => \N__39449\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39452\,
            I => \N__39446\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39449\,
            I => \N__39442\
        );

    \I__8349\ : Span4Mux_h
    port map (
            O => \N__39446\,
            I => \N__39439\
        );

    \I__8348\ : InMux
    port map (
            O => \N__39445\,
            I => \N__39436\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__39442\,
            I => \N__39433\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__39439\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__39436\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8344\ : Odrv12
    port map (
            O => \N__39433\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8343\ : InMux
    port map (
            O => \N__39426\,
            I => \bfn_16_14_0_\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39417\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39417\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__39417\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39414\,
            I => \N__39407\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39407\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39412\,
            I => \N__39404\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39401\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__39404\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8334\ : Odrv4
    port map (
            O => \N__39401\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__8333\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39390\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39390\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__39390\,
            I => \N__39386\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39383\
        );

    \I__8329\ : Span4Mux_v
    port map (
            O => \N__39386\,
            I => \N__39380\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__39383\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8327\ : Odrv4
    port map (
            O => \N__39380\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39369\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__39369\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39363\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39363\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39357\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__39357\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__8319\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39347\
        );

    \I__8318\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39347\
        );

    \I__8317\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39344\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__39347\,
            I => \N__39341\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39344\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__39341\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__39336\,
            I => \N__39332\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39326\
        );

    \I__8311\ : InMux
    port map (
            O => \N__39332\,
            I => \N__39326\
        );

    \I__8310\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39323\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__39326\,
            I => \N__39320\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__39323\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__39320\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__39312\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__39309\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__8303\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__39300\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39291\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39296\,
            I => \N__39291\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39291\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__39288\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39282\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39282\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__8293\ : InMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__8291\ : Odrv4
    port map (
            O => \N__39270\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__8290\ : InMux
    port map (
            O => \N__39267\,
            I => \N__39264\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__39264\,
            I => \N__39261\
        );

    \I__8288\ : Odrv4
    port map (
            O => \N__39261\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__8287\ : CascadeMux
    port map (
            O => \N__39258\,
            I => \N__39255\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39255\,
            I => \N__39252\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__39252\,
            I => \N__39249\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__39249\,
            I => \N__39246\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__39246\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__8282\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39240\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__8280\ : Span4Mux_h
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__39234\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__39231\,
            I => \N__39228\
        );

    \I__8277\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__39219\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39213\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__39213\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__8271\ : CascadeMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__8270\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39204\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__39204\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39201\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__39192\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39185\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39182\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39185\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__39182\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8260\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39174\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39167\
        );

    \I__8257\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39164\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__39167\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__39164\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__8253\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39153\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__39153\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__8251\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39146\
        );

    \I__8250\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39143\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39146\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39143\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8247\ : CascadeMux
    port map (
            O => \N__39138\,
            I => \N__39135\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__39132\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__8244\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39125\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39122\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39125\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__39122\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__8240\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__39114\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__8238\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__39105\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39098\
        );

    \I__8234\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39095\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__39098\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__39095\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__39090\,
            I => \N__39087\
        );

    \I__8230\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39084\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__39084\,
            I => \N__39081\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__39081\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__8227\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39074\
        );

    \I__8226\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39071\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39074\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__39071\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__39066\,
            I => \N__39063\
        );

    \I__8222\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39060\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__39060\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39054\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__39054\,
            I => \N__39051\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__39048\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__8216\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39041\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39038\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__39041\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__39038\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__39027\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__8209\ : InMux
    port map (
            O => \N__39024\,
            I => \N__39020\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__39020\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__39017\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8205\ : CascadeMux
    port map (
            O => \N__39012\,
            I => \N__39009\
        );

    \I__8204\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__39006\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__8202\ : InMux
    port map (
            O => \N__39003\,
            I => \N__38999\
        );

    \I__8201\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38996\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38999\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__38996\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38988\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38988\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__8196\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38981\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38978\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38981\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__38978\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__38973\,
            I => \N__38970\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38970\,
            I => \N__38967\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__38967\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38960\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38963\,
            I => \N__38957\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38960\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38957\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__8185\ : CascadeMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__38946\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__8180\ : Span4Mux_v
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__38934\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38927\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38930\,
            I => \N__38924\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38927\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__38924\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__38919\,
            I => \N__38916\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38913\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38907\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38904\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__38901\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38894\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38891\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__38894\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38891\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__8163\ : CascadeMux
    port map (
            O => \N__38886\,
            I => \N__38883\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38880\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38873\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38876\,
            I => \N__38870\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38873\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__38870\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8156\ : CascadeMux
    port map (
            O => \N__38865\,
            I => \N__38862\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38859\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38856\,
            I => \N__38852\
        );

    \I__8152\ : CascadeMux
    port map (
            O => \N__38855\,
            I => \N__38849\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38846\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38841\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38846\,
            I => \N__38838\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__38845\,
            I => \N__38835\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38829\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__38841\,
            I => \N__38824\
        );

    \I__8145\ : Span4Mux_v
    port map (
            O => \N__38838\,
            I => \N__38824\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38821\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38817\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38814\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38811\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38829\,
            I => \N__38808\
        );

    \I__8139\ : Sp12to4
    port map (
            O => \N__38824\,
            I => \N__38803\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38821\,
            I => \N__38803\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38800\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38817\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38814\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38811\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__38808\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8132\ : Odrv12
    port map (
            O => \N__38803\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38800\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38787\,
            I => \N__38783\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38780\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__38783\,
            I => \phase_controller_inst1.stoper_hc.N_8_0\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38780\,
            I => \phase_controller_inst1.stoper_hc.N_8_0\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38767\
        );

    \I__8125\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38764\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38761\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38754\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38754\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38770\,
            I => \N__38754\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38767\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38764\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38761\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38754\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__8116\ : IoInMux
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__8114\ : IoSpan4Mux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__8113\ : Span4Mux_s2_v
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__8112\ : Sp12to4
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__8111\ : Span12Mux_v
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__8110\ : Span12Mux_v
    port map (
            O => \N__38727\,
            I => \N__38723\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38720\
        );

    \I__8108\ : Odrv12
    port map (
            O => \N__38723\,
            I => test22_c
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38720\,
            I => test22_c
        );

    \I__8106\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38711\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38708\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__38711\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__38708\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38703\,
            I => \N__38699\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38696\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38699\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38696\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__38682\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__8094\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38675\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38671\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38675\,
            I => \N__38668\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38665\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38671\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8089\ : Odrv12
    port map (
            O => \N__38668\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38665\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__8087\ : IoInMux
    port map (
            O => \N__38658\,
            I => \N__38655\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__38655\,
            I => \N__38652\
        );

    \I__8085\ : Span4Mux_s3_v
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__8083\ : Span4Mux_v
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__38643\,
            I => \current_shift_inst.timer_s1.N_339_i\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__38640\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__38634\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__38631\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38625\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38625\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__38619\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38609\
        );

    \I__8071\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38606\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__38609\,
            I => \N__38603\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38606\,
            I => \N__38599\
        );

    \I__8068\ : Span4Mux_v
    port map (
            O => \N__38603\,
            I => \N__38596\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38602\,
            I => \N__38593\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__38599\,
            I => \N__38589\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__38596\,
            I => \N__38586\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__38593\,
            I => \N__38583\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38580\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__38589\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__38586\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8060\ : Odrv4
    port map (
            O => \N__38583\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38580\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38566\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38563\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38560\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__38566\,
            I => \N__38555\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__38563\,
            I => \N__38555\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__38560\,
            I => \N__38552\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__38555\,
            I => \N__38547\
        );

    \I__8051\ : Span4Mux_h
    port map (
            O => \N__38552\,
            I => \N__38547\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__38547\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__38544\,
            I => \N__38541\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__8046\ : Odrv12
    port map (
            O => \N__38535\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38510\
        );

    \I__8044\ : InMux
    port map (
            O => \N__38531\,
            I => \N__38510\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38530\,
            I => \N__38510\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38501\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38501\
        );

    \I__8040\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38501\
        );

    \I__8039\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38501\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38494\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38491\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38486\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38486\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38483\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38478\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38478\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38475\
        );

    \I__8030\ : InMux
    port map (
            O => \N__38517\,
            I => \N__38472\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__38510\,
            I => \N__38467\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__38501\,
            I => \N__38467\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38462\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38462\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38457\
        );

    \I__8024\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38457\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__38494\,
            I => \N__38452\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38491\,
            I => \N__38452\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38486\,
            I => \N__38449\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__38483\,
            I => \N__38440\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38478\,
            I => \N__38440\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__38475\,
            I => \N__38440\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38472\,
            I => \N__38433\
        );

    \I__8016\ : Span4Mux_v
    port map (
            O => \N__38467\,
            I => \N__38433\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38462\,
            I => \N__38433\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__38457\,
            I => \N__38423\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__38452\,
            I => \N__38423\
        );

    \I__8012\ : Span4Mux_v
    port map (
            O => \N__38449\,
            I => \N__38423\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38418\
        );

    \I__8010\ : InMux
    port map (
            O => \N__38447\,
            I => \N__38418\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__38440\,
            I => \N__38413\
        );

    \I__8008\ : Span4Mux_v
    port map (
            O => \N__38433\,
            I => \N__38413\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38410\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38405\
        );

    \I__8005\ : InMux
    port map (
            O => \N__38430\,
            I => \N__38405\
        );

    \I__8004\ : Odrv4
    port map (
            O => \N__38423\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38418\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__38413\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38410\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38405\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__38394\,
            I => \N__38391\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38388\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__38388\,
            I => \N__38384\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38381\
        );

    \I__7995\ : Span4Mux_h
    port map (
            O => \N__38384\,
            I => \N__38378\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38381\,
            I => \N__38373\
        );

    \I__7993\ : Span4Mux_h
    port map (
            O => \N__38378\,
            I => \N__38370\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38367\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38376\,
            I => \N__38364\
        );

    \I__7990\ : Odrv12
    port map (
            O => \N__38373\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__38370\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__38367\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__38364\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__7986\ : CascadeMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__7985\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38348\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38351\,
            I => \N__38344\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38348\,
            I => \N__38341\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38338\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38344\,
            I => \N__38335\
        );

    \I__7980\ : Span4Mux_h
    port map (
            O => \N__38341\,
            I => \N__38332\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__38338\,
            I => \N__38329\
        );

    \I__7978\ : Span4Mux_h
    port map (
            O => \N__38335\,
            I => \N__38326\
        );

    \I__7977\ : Odrv4
    port map (
            O => \N__38332\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7976\ : Odrv12
    port map (
            O => \N__38329\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__38326\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38313\
        );

    \I__7972\ : Span4Mux_v
    port map (
            O => \N__38313\,
            I => \N__38310\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__38310\,
            I => \N__38307\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__38307\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__7969\ : InMux
    port map (
            O => \N__38304\,
            I => \N__38300\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38297\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__38300\,
            I => \N__38291\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__38297\,
            I => \N__38291\
        );

    \I__7965\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38288\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__38291\,
            I => \N__38283\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__38288\,
            I => \N__38283\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__38283\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38276\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38273\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__38276\,
            I => \N__38266\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__38273\,
            I => \N__38266\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38261\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38261\
        );

    \I__7955\ : Span4Mux_v
    port map (
            O => \N__38266\,
            I => \N__38258\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__38261\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__38258\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7952\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38245\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38252\,
            I => \N__38245\
        );

    \I__7950\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38242\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38239\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38236\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38242\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__38239\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7945\ : Odrv12
    port map (
            O => \N__38236\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38229\,
            I => \N__38226\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__7942\ : Span4Mux_s3_h
    port map (
            O => \N__38223\,
            I => \N__38219\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38216\
        );

    \I__7940\ : Sp12to4
    port map (
            O => \N__38219\,
            I => \N__38213\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38216\,
            I => \N__38210\
        );

    \I__7938\ : Span12Mux_s11_v
    port map (
            O => \N__38213\,
            I => \N__38207\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__38210\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__7936\ : Odrv12
    port map (
            O => \N__38207\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__7935\ : InMux
    port map (
            O => \N__38202\,
            I => \N__38199\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38199\,
            I => \N__38196\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__7932\ : Sp12to4
    port map (
            O => \N__38193\,
            I => \N__38190\
        );

    \I__7931\ : Odrv12
    port map (
            O => \N__38190\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38182\
        );

    \I__7929\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38179\
        );

    \I__7928\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38175\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38182\,
            I => \N__38170\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__38179\,
            I => \N__38170\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38167\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38175\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7923\ : Odrv4
    port map (
            O => \N__38170\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__38167\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7921\ : CEMux
    port map (
            O => \N__38160\,
            I => \N__38157\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__38154\,
            I => \N__38150\
        );

    \I__7918\ : InMux
    port map (
            O => \N__38153\,
            I => \N__38147\
        );

    \I__7917\ : Sp12to4
    port map (
            O => \N__38150\,
            I => \N__38142\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38142\
        );

    \I__7915\ : Span12Mux_v
    port map (
            O => \N__38142\,
            I => \N__38139\
        );

    \I__7914\ : Odrv12
    port map (
            O => \N__38139\,
            I => \S1_RNI9RLH\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__38136\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__7912\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__7910\ : Span4Mux_h
    port map (
            O => \N__38127\,
            I => \N__38124\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__38124\,
            I => \current_shift_inst.PI_CTRL.N_286\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38118\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__7906\ : Odrv12
    port map (
            O => \N__38115\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38108\
        );

    \I__7904\ : InMux
    port map (
            O => \N__38111\,
            I => \N__38105\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__38108\,
            I => \N__38102\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__38105\,
            I => \N__38098\
        );

    \I__7901\ : Span4Mux_h
    port map (
            O => \N__38102\,
            I => \N__38095\
        );

    \I__7900\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38092\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__38098\,
            I => \N__38085\
        );

    \I__7898\ : Span4Mux_v
    port map (
            O => \N__38095\,
            I => \N__38085\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__38092\,
            I => \N__38085\
        );

    \I__7896\ : Span4Mux_h
    port map (
            O => \N__38085\,
            I => \N__38081\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38078\
        );

    \I__7894\ : Odrv4
    port map (
            O => \N__38081\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__38078\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38073\,
            I => \N__38070\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__38070\,
            I => \N__38067\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__38067\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__7889\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38061\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__38057\
        );

    \I__7887\ : InMux
    port map (
            O => \N__38060\,
            I => \N__38054\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__38057\,
            I => \N__38049\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__38054\,
            I => \N__38049\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__38049\,
            I => \N__38044\
        );

    \I__7883\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38041\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38038\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__38044\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__38041\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__38038\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__7878\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38026\
        );

    \I__7877\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38023\
        );

    \I__7876\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38020\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38017\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__38014\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__38020\,
            I => \N__38011\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__38017\,
            I => \N__38008\
        );

    \I__7871\ : Span4Mux_h
    port map (
            O => \N__38014\,
            I => \N__38005\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__38011\,
            I => \N__38002\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__38008\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__38005\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__38002\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37992\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37992\,
            I => \N__37989\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__37989\,
            I => \N__37986\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__37986\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__7862\ : CascadeMux
    port map (
            O => \N__37983\,
            I => \N__37979\
        );

    \I__7861\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37976\
        );

    \I__7860\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37973\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__37976\,
            I => \N__37970\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__37973\,
            I => \N__37967\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__37970\,
            I => \N__37962\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__37967\,
            I => \N__37962\
        );

    \I__7855\ : Span4Mux_h
    port map (
            O => \N__37962\,
            I => \N__37957\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37954\
        );

    \I__7853\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37951\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__37957\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37954\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37951\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37941\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37941\,
            I => \N__37937\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37934\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__37937\,
            I => \N__37930\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37934\,
            I => \N__37927\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37924\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__37930\,
            I => \N__37921\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__37927\,
            I => \N__37918\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37924\,
            I => \N__37915\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__37921\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__37918\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7838\ : Odrv4
    port map (
            O => \N__37915\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37902\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37899\
        );

    \I__7834\ : Span4Mux_h
    port map (
            O => \N__37899\,
            I => \N__37896\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__37896\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__37893\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37890\,
            I => \N__37884\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37884\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37884\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37874\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37874\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37871\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37874\,
            I => \N__37868\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__37871\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__37868\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__37863\,
            I => \N__37859\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37853\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37853\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37850\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__37853\,
            I => \N__37847\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37850\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__37847\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__37842\,
            I => \N__37838\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37833\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37833\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__37833\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__7811\ : CascadeMux
    port map (
            O => \N__37830\,
            I => \N__37827\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37827\,
            I => \N__37823\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__37826\,
            I => \N__37820\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37817\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37814\
        );

    \I__7806\ : Span4Mux_h
    port map (
            O => \N__37817\,
            I => \N__37811\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37808\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__37811\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__37808\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37803\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37800\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37797\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37794\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37786\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37781\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37781\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37786\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__37781\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__37776\,
            I => \N__37771\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37768\
        );

    \I__7791\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37763\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37763\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37768\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37763\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7787\ : CascadeMux
    port map (
            O => \N__37758\,
            I => \N__37755\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37755\,
            I => \N__37749\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37749\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37749\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37740\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37740\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37740\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37737\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7779\ : InMux
    port map (
            O => \N__37734\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37731\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37728\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37725\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37717\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37714\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37711\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37708\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37714\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37711\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7769\ : Odrv4
    port map (
            O => \N__37708\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37701\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37693\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37690\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37687\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37693\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__37690\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37687\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37680\,
            I => \bfn_15_8_0_\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37677\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37674\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37671\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37668\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37665\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37662\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37659\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37656\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37653\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37650\,
            I => \bfn_15_7_0_\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37647\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37644\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__37641\,
            I => \N__37637\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__37640\,
            I => \N__37634\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37629\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37629\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37629\,
            I => \phase_controller_inst1.stoper_hc.N_45_i\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37626\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37623\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37620\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__7740\ : InMux
    port map (
            O => \N__37617\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37614\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__7738\ : InMux
    port map (
            O => \N__37611\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37608\,
            I => \bfn_15_6_0_\
        );

    \I__7736\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37602\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__37602\,
            I => \phase_controller_inst1.stoper_hc.N_27\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37596\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__37590\,
            I => \N__37587\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__37587\,
            I => il_max_comp1_c
        );

    \I__7729\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37581\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__37581\,
            I => \N__37576\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37569\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37569\
        );

    \I__7725\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37566\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37575\,
            I => \N__37563\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37574\,
            I => \N__37560\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__37569\,
            I => \phase_controller_inst1.N_175_1\
        );

    \I__7721\ : Odrv4
    port map (
            O => \N__37566\,
            I => \phase_controller_inst1.N_175_1\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__37563\,
            I => \phase_controller_inst1.N_175_1\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37560\,
            I => \phase_controller_inst1.N_175_1\
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__37551\,
            I => \phase_controller_inst1.stoper_hc.N_8_0_cascade_\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37545\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37545\,
            I => \phase_controller_inst1.stoper_hc.m12_ns_1\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37542\,
            I => \N__37535\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37535\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37530\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37527\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37524\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37533\,
            I => \N__37521\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__37530\,
            I => \N__37518\
        );

    \I__7708\ : Span4Mux_h
    port map (
            O => \N__37527\,
            I => \N__37515\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37524\,
            I => \N__37510\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__37521\,
            I => \N__37510\
        );

    \I__7705\ : Span12Mux_h
    port map (
            O => \N__37518\,
            I => \N__37507\
        );

    \I__7704\ : IoSpan4Mux
    port map (
            O => \N__37515\,
            I => \N__37502\
        );

    \I__7703\ : IoSpan4Mux
    port map (
            O => \N__37510\,
            I => \N__37502\
        );

    \I__7702\ : Odrv12
    port map (
            O => \N__37507\,
            I => il_min_comp1_c
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__37502\,
            I => il_min_comp1_c
        );

    \I__7700\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37494\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37494\,
            I => \phase_controller_inst1.N_14_0\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__7697\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37485\,
            I => \N__37482\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__37482\,
            I => \phase_controller_inst1.N_13_0\
        );

    \I__7694\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37476\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37473\
        );

    \I__7692\ : Span4Mux_v
    port map (
            O => \N__37473\,
            I => \N__37467\
        );

    \I__7691\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37464\
        );

    \I__7690\ : CascadeMux
    port map (
            O => \N__37471\,
            I => \N__37459\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37456\
        );

    \I__7688\ : Sp12to4
    port map (
            O => \N__37467\,
            I => \N__37453\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__37464\,
            I => \N__37450\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37447\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37442\
        );

    \I__7684\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37442\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37437\
        );

    \I__7682\ : Span12Mux_v
    port map (
            O => \N__37453\,
            I => \N__37437\
        );

    \I__7681\ : Span4Mux_h
    port map (
            O => \N__37450\,
            I => \N__37434\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__37447\,
            I => \N__37431\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37442\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7678\ : Odrv12
    port map (
            O => \N__37437\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7677\ : Odrv4
    port map (
            O => \N__37434\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__37431\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37419\,
            I => \phase_controller_inst2.m21\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37412\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__37415\,
            I => \N__37409\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__37412\,
            I => \N__37406\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37403\
        );

    \I__7669\ : Sp12to4
    port map (
            O => \N__37406\,
            I => \N__37398\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37395\
        );

    \I__7667\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37392\
        );

    \I__7666\ : CascadeMux
    port map (
            O => \N__37401\,
            I => \N__37389\
        );

    \I__7665\ : Span12Mux_s8_v
    port map (
            O => \N__37398\,
            I => \N__37384\
        );

    \I__7664\ : Span4Mux_v
    port map (
            O => \N__37395\,
            I => \N__37379\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__37392\,
            I => \N__37379\
        );

    \I__7662\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37376\
        );

    \I__7661\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37373\
        );

    \I__7660\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37370\
        );

    \I__7659\ : Span12Mux_v
    port map (
            O => \N__37384\,
            I => \N__37367\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__37379\,
            I => \N__37364\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__37376\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__37373\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__37370\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7654\ : Odrv12
    port map (
            O => \N__37367\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__37364\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__37350\,
            I => \phase_controller_inst2.time_passed_er_RNI23UO1\
        );

    \I__7650\ : IoInMux
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__37344\,
            I => \N__37341\
        );

    \I__7648\ : Span4Mux_s2_v
    port map (
            O => \N__37341\,
            I => \N__37338\
        );

    \I__7647\ : Sp12to4
    port map (
            O => \N__37338\,
            I => \N__37335\
        );

    \I__7646\ : Span12Mux_h
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__7645\ : Span12Mux_v
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__7644\ : Span12Mux_v
    port map (
            O => \N__37329\,
            I => \N__37325\
        );

    \I__7643\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37322\
        );

    \I__7642\ : Odrv12
    port map (
            O => \N__37325\,
            I => s1_phy_c
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37322\,
            I => s1_phy_c
        );

    \I__7640\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37313\
        );

    \I__7639\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37310\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37307\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__37310\,
            I => \N__37304\
        );

    \I__7636\ : Span4Mux_v
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__37304\,
            I => \N__37298\
        );

    \I__7634\ : Sp12to4
    port map (
            O => \N__37301\,
            I => \N__37295\
        );

    \I__7633\ : Span4Mux_h
    port map (
            O => \N__37298\,
            I => \N__37292\
        );

    \I__7632\ : Span12Mux_h
    port map (
            O => \N__37295\,
            I => \N__37289\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__37292\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__7630\ : Odrv12
    port map (
            O => \N__37289\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37284\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__37278\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__7626\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37271\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37268\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__37271\,
            I => \N__37265\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__37268\,
            I => \N__37262\
        );

    \I__7622\ : Span4Mux_v
    port map (
            O => \N__37265\,
            I => \N__37259\
        );

    \I__7621\ : Span4Mux_s3_h
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__7620\ : Sp12to4
    port map (
            O => \N__37259\,
            I => \N__37253\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__37256\,
            I => \N__37250\
        );

    \I__7618\ : Span12Mux_s7_h
    port map (
            O => \N__37253\,
            I => \N__37245\
        );

    \I__7617\ : Sp12to4
    port map (
            O => \N__37250\,
            I => \N__37245\
        );

    \I__7616\ : Span12Mux_v
    port map (
            O => \N__37245\,
            I => \N__37242\
        );

    \I__7615\ : Odrv12
    port map (
            O => \N__37242\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__7614\ : InMux
    port map (
            O => \N__37239\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__7613\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37233\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__37233\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__7611\ : InMux
    port map (
            O => \N__37230\,
            I => \N__37227\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37227\,
            I => \N__37223\
        );

    \I__7609\ : InMux
    port map (
            O => \N__37226\,
            I => \N__37220\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__37223\,
            I => \N__37217\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__37220\,
            I => \N__37214\
        );

    \I__7606\ : Sp12to4
    port map (
            O => \N__37217\,
            I => \N__37211\
        );

    \I__7605\ : Span4Mux_v
    port map (
            O => \N__37214\,
            I => \N__37208\
        );

    \I__7604\ : Span12Mux_s6_h
    port map (
            O => \N__37211\,
            I => \N__37205\
        );

    \I__7603\ : Sp12to4
    port map (
            O => \N__37208\,
            I => \N__37200\
        );

    \I__7602\ : Span12Mux_v
    port map (
            O => \N__37205\,
            I => \N__37200\
        );

    \I__7601\ : Odrv12
    port map (
            O => \N__37200\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37197\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__7599\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37191\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__37191\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__7597\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37185\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__37185\,
            I => \N__37181\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37178\
        );

    \I__7594\ : Sp12to4
    port map (
            O => \N__37181\,
            I => \N__37175\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37172\
        );

    \I__7592\ : Span12Mux_v
    port map (
            O => \N__37175\,
            I => \N__37169\
        );

    \I__7591\ : Span12Mux_v
    port map (
            O => \N__37172\,
            I => \N__37166\
        );

    \I__7590\ : Span12Mux_h
    port map (
            O => \N__37169\,
            I => \N__37163\
        );

    \I__7589\ : Odrv12
    port map (
            O => \N__37166\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7588\ : Odrv12
    port map (
            O => \N__37163\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37158\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37155\,
            I => \N__37152\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__37152\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__7584\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37145\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37142\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37139\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37136\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__37139\,
            I => \N__37133\
        );

    \I__7579\ : Span12Mux_v
    port map (
            O => \N__37136\,
            I => \N__37130\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__37133\,
            I => \N__37127\
        );

    \I__7577\ : Span12Mux_h
    port map (
            O => \N__37130\,
            I => \N__37124\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__37127\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__7575\ : Odrv12
    port map (
            O => \N__37124\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37119\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37112\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37109\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37112\,
            I => \current_shift_inst.control_input_31\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37109\,
            I => \current_shift_inst.control_input_31\
        );

    \I__7569\ : InMux
    port map (
            O => \N__37104\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37101\,
            I => \N__37098\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__37098\,
            I => \N__37095\
        );

    \I__7566\ : Span4Mux_h
    port map (
            O => \N__37095\,
            I => \N__37092\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__37089\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__7563\ : IoInMux
    port map (
            O => \N__37086\,
            I => \N__37083\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__37083\,
            I => \N__37080\
        );

    \I__7561\ : Span12Mux_s5_v
    port map (
            O => \N__37080\,
            I => \N__37077\
        );

    \I__7560\ : Odrv12
    port map (
            O => \N__37077\,
            I => s2_phy_c
        );

    \I__7559\ : InMux
    port map (
            O => \N__37074\,
            I => \N__37071\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__37071\,
            I => \N__37068\
        );

    \I__7557\ : Odrv4
    port map (
            O => \N__37068\,
            I => \phase_controller_inst1.stoper_hc.m19_ns_1\
        );

    \I__7556\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37062\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__37062\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37059\,
            I => \N__37056\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__7552\ : Span4Mux_s2_h
    port map (
            O => \N__37053\,
            I => \N__37049\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37046\
        );

    \I__7550\ : Sp12to4
    port map (
            O => \N__37049\,
            I => \N__37043\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37038\
        );

    \I__7548\ : Span12Mux_v
    port map (
            O => \N__37043\,
            I => \N__37038\
        );

    \I__7547\ : Span12Mux_h
    port map (
            O => \N__37038\,
            I => \N__37035\
        );

    \I__7546\ : Odrv12
    port map (
            O => \N__37035\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__7545\ : InMux
    port map (
            O => \N__37032\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__7544\ : InMux
    port map (
            O => \N__37029\,
            I => \N__37026\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__37026\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37023\,
            I => \N__37019\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37022\,
            I => \N__37016\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37019\,
            I => \N__37013\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37010\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__37013\,
            I => \N__37007\
        );

    \I__7537\ : Span12Mux_s2_h
    port map (
            O => \N__37010\,
            I => \N__37004\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__37007\,
            I => \N__37001\
        );

    \I__7535\ : Span12Mux_h
    port map (
            O => \N__37004\,
            I => \N__36998\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__37001\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7533\ : Odrv12
    port map (
            O => \N__36998\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36993\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36987\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__36987\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36980\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36974\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36971\
        );

    \I__7525\ : Sp12to4
    port map (
            O => \N__36974\,
            I => \N__36968\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__36971\,
            I => \N__36965\
        );

    \I__7523\ : Span12Mux_v
    port map (
            O => \N__36968\,
            I => \N__36962\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__36965\,
            I => \N__36959\
        );

    \I__7521\ : Span12Mux_h
    port map (
            O => \N__36962\,
            I => \N__36956\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__36959\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__7519\ : Odrv12
    port map (
            O => \N__36956\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36951\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__36945\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36939\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36939\,
            I => \N__36935\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36932\
        );

    \I__7512\ : Span4Mux_v
    port map (
            O => \N__36935\,
            I => \N__36929\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36926\
        );

    \I__7510\ : Sp12to4
    port map (
            O => \N__36929\,
            I => \N__36921\
        );

    \I__7509\ : Span12Mux_v
    port map (
            O => \N__36926\,
            I => \N__36921\
        );

    \I__7508\ : Span12Mux_h
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__7507\ : Odrv12
    port map (
            O => \N__36918\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36915\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36909\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__36909\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36903\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36900\
        );

    \I__7501\ : Span4Mux_s3_h
    port map (
            O => \N__36900\,
            I => \N__36896\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36893\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__36896\,
            I => \N__36890\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36893\,
            I => \N__36885\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__36890\,
            I => \N__36885\
        );

    \I__7496\ : Sp12to4
    port map (
            O => \N__36885\,
            I => \N__36882\
        );

    \I__7495\ : Odrv12
    port map (
            O => \N__36882\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36879\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36873\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36873\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36866\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36863\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__36866\,
            I => \N__36860\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36863\,
            I => \N__36857\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__36860\,
            I => \N__36854\
        );

    \I__7486\ : Span4Mux_h
    port map (
            O => \N__36857\,
            I => \N__36851\
        );

    \I__7485\ : Span4Mux_s1_h
    port map (
            O => \N__36854\,
            I => \N__36848\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__36851\,
            I => \N__36845\
        );

    \I__7483\ : Sp12to4
    port map (
            O => \N__36848\,
            I => \N__36842\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__36845\,
            I => \N__36839\
        );

    \I__7481\ : Span12Mux_h
    port map (
            O => \N__36842\,
            I => \N__36836\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__36839\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__7479\ : Odrv12
    port map (
            O => \N__36836\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36831\,
            I => \bfn_14_21_0_\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36825\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36825\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36818\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36815\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36818\,
            I => \N__36812\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__36815\,
            I => \N__36809\
        );

    \I__7471\ : Span4Mux_v
    port map (
            O => \N__36812\,
            I => \N__36806\
        );

    \I__7470\ : Span4Mux_v
    port map (
            O => \N__36809\,
            I => \N__36803\
        );

    \I__7469\ : Sp12to4
    port map (
            O => \N__36806\,
            I => \N__36800\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__36803\,
            I => \N__36797\
        );

    \I__7467\ : Span12Mux_s2_h
    port map (
            O => \N__36800\,
            I => \N__36794\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__36797\,
            I => \N__36791\
        );

    \I__7465\ : Span12Mux_h
    port map (
            O => \N__36794\,
            I => \N__36788\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__36791\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__7463\ : Odrv12
    port map (
            O => \N__36788\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36783\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36777\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36771\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36771\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36768\,
            I => \N__36765\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36765\,
            I => \N__36762\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__36762\,
            I => \N__36758\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36755\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__36758\,
            I => \N__36752\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36749\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__36752\,
            I => \N__36746\
        );

    \I__7450\ : Span12Mux_s11_v
    port map (
            O => \N__36749\,
            I => \N__36743\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__36746\,
            I => \N__36740\
        );

    \I__7448\ : Odrv12
    port map (
            O => \N__36743\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__36740\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36735\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36729\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36729\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36722\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36719\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36716\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__36719\,
            I => \N__36713\
        );

    \I__7439\ : Span4Mux_v
    port map (
            O => \N__36716\,
            I => \N__36710\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__36713\,
            I => \N__36707\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__36710\,
            I => \N__36704\
        );

    \I__7436\ : Span4Mux_h
    port map (
            O => \N__36707\,
            I => \N__36701\
        );

    \I__7435\ : Sp12to4
    port map (
            O => \N__36704\,
            I => \N__36698\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__36701\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7433\ : Odrv12
    port map (
            O => \N__36698\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36693\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36687\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36687\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36681\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36677\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36674\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__36677\,
            I => \N__36671\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36668\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__36671\,
            I => \N__36665\
        );

    \I__7423\ : Span12Mux_s11_v
    port map (
            O => \N__36668\,
            I => \N__36662\
        );

    \I__7422\ : Odrv4
    port map (
            O => \N__36665\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7421\ : Odrv12
    port map (
            O => \N__36662\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36657\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36651\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36651\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36645\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__36645\,
            I => \N__36641\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36644\,
            I => \N__36638\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36635\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36638\,
            I => \N__36632\
        );

    \I__7412\ : Span4Mux_h
    port map (
            O => \N__36635\,
            I => \N__36629\
        );

    \I__7411\ : Span12Mux_s11_h
    port map (
            O => \N__36632\,
            I => \N__36626\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__36629\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7409\ : Odrv12
    port map (
            O => \N__36626\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36621\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36615\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36615\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36609\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36606\
        );

    \I__7403\ : Span4Mux_s3_h
    port map (
            O => \N__36606\,
            I => \N__36602\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36599\
        );

    \I__7401\ : Sp12to4
    port map (
            O => \N__36602\,
            I => \N__36596\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36591\
        );

    \I__7399\ : Span12Mux_v
    port map (
            O => \N__36596\,
            I => \N__36591\
        );

    \I__7398\ : Odrv12
    port map (
            O => \N__36591\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36588\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36585\,
            I => \N__36582\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36582\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36575\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36578\,
            I => \N__36572\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__36575\,
            I => \N__36569\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__36572\,
            I => \N__36566\
        );

    \I__7390\ : Span4Mux_v
    port map (
            O => \N__36569\,
            I => \N__36563\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__36566\,
            I => \N__36560\
        );

    \I__7388\ : Sp12to4
    port map (
            O => \N__36563\,
            I => \N__36557\
        );

    \I__7387\ : Span4Mux_h
    port map (
            O => \N__36560\,
            I => \N__36554\
        );

    \I__7386\ : Span12Mux_s10_h
    port map (
            O => \N__36557\,
            I => \N__36551\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__36554\,
            I => \N__36548\
        );

    \I__7384\ : Span12Mux_v
    port map (
            O => \N__36551\,
            I => \N__36545\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__36548\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7382\ : Odrv12
    port map (
            O => \N__36545\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36540\,
            I => \bfn_14_20_0_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36534\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36534\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36528\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__36528\,
            I => \N__36525\
        );

    \I__7376\ : Span4Mux_s2_h
    port map (
            O => \N__36525\,
            I => \N__36521\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36518\
        );

    \I__7374\ : Sp12to4
    port map (
            O => \N__36521\,
            I => \N__36515\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36510\
        );

    \I__7372\ : Span12Mux_v
    port map (
            O => \N__36515\,
            I => \N__36510\
        );

    \I__7371\ : Span12Mux_h
    port map (
            O => \N__36510\,
            I => \N__36507\
        );

    \I__7370\ : Odrv12
    port map (
            O => \N__36507\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36504\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__7368\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36498\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__36498\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36491\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36488\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__36491\,
            I => \N__36485\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__36488\,
            I => \N__36482\
        );

    \I__7362\ : Span4Mux_h
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__7361\ : Span4Mux_v
    port map (
            O => \N__36482\,
            I => \N__36476\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__36479\,
            I => \N__36473\
        );

    \I__7359\ : Sp12to4
    port map (
            O => \N__36476\,
            I => \N__36470\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__36473\,
            I => \N__36467\
        );

    \I__7357\ : Span12Mux_h
    port map (
            O => \N__36470\,
            I => \N__36464\
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__36467\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__36464\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36459\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36453\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__36453\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36447\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36444\
        );

    \I__7349\ : Span4Mux_s2_h
    port map (
            O => \N__36444\,
            I => \N__36440\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36437\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__36440\,
            I => \N__36434\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__36437\,
            I => \N__36431\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__36434\,
            I => \N__36428\
        );

    \I__7344\ : Span12Mux_v
    port map (
            O => \N__36431\,
            I => \N__36425\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__36428\,
            I => \N__36422\
        );

    \I__7342\ : Odrv12
    port map (
            O => \N__36425\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__7341\ : Odrv4
    port map (
            O => \N__36422\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__7340\ : InMux
    port map (
            O => \N__36417\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36411\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__36411\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36408\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36402\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__36402\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36396\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36396\,
            I => \N__36392\
        );

    \I__7332\ : InMux
    port map (
            O => \N__36395\,
            I => \N__36389\
        );

    \I__7331\ : Span4Mux_h
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__36386\,
            I => \N__36380\
        );

    \I__7328\ : Span12Mux_v
    port map (
            O => \N__36383\,
            I => \N__36377\
        );

    \I__7327\ : Odrv4
    port map (
            O => \N__36380\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__7326\ : Odrv12
    port map (
            O => \N__36377\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36372\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__7324\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36366\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36366\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36359\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36353\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36356\,
            I => \N__36350\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__36353\,
            I => \N__36347\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__36350\,
            I => \N__36344\
        );

    \I__7316\ : Span4Mux_v
    port map (
            O => \N__36347\,
            I => \N__36341\
        );

    \I__7315\ : Span4Mux_h
    port map (
            O => \N__36344\,
            I => \N__36338\
        );

    \I__7314\ : Sp12to4
    port map (
            O => \N__36341\,
            I => \N__36335\
        );

    \I__7313\ : Odrv4
    port map (
            O => \N__36338\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7312\ : Odrv12
    port map (
            O => \N__36335\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36330\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36324\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36324\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36317\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36314\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__36317\,
            I => \N__36311\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__36314\,
            I => \N__36308\
        );

    \I__7304\ : Span12Mux_s11_h
    port map (
            O => \N__36311\,
            I => \N__36305\
        );

    \I__7303\ : Odrv12
    port map (
            O => \N__36308\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__7302\ : Odrv12
    port map (
            O => \N__36305\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36300\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__7300\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__36294\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36291\,
            I => \bfn_14_19_0_\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36285\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36285\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36282\,
            I => \N__36279\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__7293\ : Span4Mux_s2_h
    port map (
            O => \N__36276\,
            I => \N__36272\
        );

    \I__7292\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36269\
        );

    \I__7291\ : Span4Mux_h
    port map (
            O => \N__36272\,
            I => \N__36266\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__36269\,
            I => \N__36263\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__36266\,
            I => \N__36260\
        );

    \I__7288\ : Span12Mux_s9_h
    port map (
            O => \N__36263\,
            I => \N__36257\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__36260\,
            I => \N__36254\
        );

    \I__7286\ : Odrv12
    port map (
            O => \N__36257\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__36254\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36249\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36243\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__36243\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36240\,
            I => \N__36237\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__7279\ : Span4Mux_s3_h
    port map (
            O => \N__36234\,
            I => \N__36230\
        );

    \I__7278\ : InMux
    port map (
            O => \N__36233\,
            I => \N__36227\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__36230\,
            I => \N__36224\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__36227\,
            I => \N__36221\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__36224\,
            I => \N__36218\
        );

    \I__7274\ : Span12Mux_s8_h
    port map (
            O => \N__36221\,
            I => \N__36215\
        );

    \I__7273\ : Sp12to4
    port map (
            O => \N__36218\,
            I => \N__36212\
        );

    \I__7272\ : Odrv12
    port map (
            O => \N__36215\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7271\ : Odrv12
    port map (
            O => \N__36212\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36207\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__7269\ : InMux
    port map (
            O => \N__36204\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__7268\ : InMux
    port map (
            O => \N__36201\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__7267\ : CEMux
    port map (
            O => \N__36198\,
            I => \N__36174\
        );

    \I__7266\ : CEMux
    port map (
            O => \N__36197\,
            I => \N__36174\
        );

    \I__7265\ : CEMux
    port map (
            O => \N__36196\,
            I => \N__36174\
        );

    \I__7264\ : CEMux
    port map (
            O => \N__36195\,
            I => \N__36174\
        );

    \I__7263\ : CEMux
    port map (
            O => \N__36194\,
            I => \N__36174\
        );

    \I__7262\ : CEMux
    port map (
            O => \N__36193\,
            I => \N__36174\
        );

    \I__7261\ : CEMux
    port map (
            O => \N__36192\,
            I => \N__36174\
        );

    \I__7260\ : CEMux
    port map (
            O => \N__36191\,
            I => \N__36174\
        );

    \I__7259\ : GlobalMux
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__7258\ : gio2CtrlBuf
    port map (
            O => \N__36171\,
            I => \current_shift_inst.timer_s1.N_339_i_g\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36168\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36161\
        );

    \I__7255\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36157\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__36161\,
            I => \N__36154\
        );

    \I__7253\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36151\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__36148\
        );

    \I__7251\ : Span4Mux_h
    port map (
            O => \N__36154\,
            I => \N__36145\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36142\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__36148\,
            I => \N__36139\
        );

    \I__7248\ : Span4Mux_h
    port map (
            O => \N__36145\,
            I => \N__36134\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__36142\,
            I => \N__36134\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__36139\,
            I => \N__36131\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__36134\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__36131\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__7243\ : CascadeMux
    port map (
            O => \N__36126\,
            I => \N__36122\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36118\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36115\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36112\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__36109\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36104\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__36112\,
            I => \N__36104\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__36109\,
            I => \N__36098\
        );

    \I__7235\ : Span4Mux_h
    port map (
            O => \N__36104\,
            I => \N__36098\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36095\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__36098\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__36095\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__7231\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__7229\ : Span4Mux_h
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__36081\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__7227\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36074\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36077\,
            I => \N__36071\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__36068\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36062\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__36068\,
            I => \N__36062\
        );

    \I__7222\ : InMux
    port map (
            O => \N__36067\,
            I => \N__36059\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__36062\,
            I => \N__36053\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__36053\
        );

    \I__7219\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36050\
        );

    \I__7218\ : Odrv4
    port map (
            O => \N__36053\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__36050\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__7216\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36042\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__36042\,
            I => \N__36039\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__36039\,
            I => \N__36036\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__36036\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__7212\ : InMux
    port map (
            O => \N__36033\,
            I => \N__36030\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__36030\,
            I => \current_shift_inst.control_input_1\
        );

    \I__7210\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36024\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__36024\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__7208\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36018\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__36018\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__7206\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36011\
        );

    \I__7205\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36008\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__36011\,
            I => \N__36005\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__36002\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__36005\,
            I => \N__35999\
        );

    \I__7201\ : Span4Mux_v
    port map (
            O => \N__36002\,
            I => \N__35996\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__35999\,
            I => \N__35993\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__7198\ : Span4Mux_h
    port map (
            O => \N__35993\,
            I => \N__35987\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__35990\,
            I => \N__35982\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__35987\,
            I => \N__35982\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__35982\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35979\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35973\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35973\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35967\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35963\
        );

    \I__7189\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35960\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__35963\,
            I => \N__35957\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__35960\,
            I => \N__35954\
        );

    \I__7186\ : Sp12to4
    port map (
            O => \N__35957\,
            I => \N__35951\
        );

    \I__7185\ : Span4Mux_h
    port map (
            O => \N__35954\,
            I => \N__35948\
        );

    \I__7184\ : Span12Mux_s11_h
    port map (
            O => \N__35951\,
            I => \N__35945\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__35948\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__7182\ : Odrv12
    port map (
            O => \N__35945\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35940\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__35937\,
            I => \N__35933\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__35936\,
            I => \N__35930\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35927\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35924\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35921\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35918\
        );

    \I__7174\ : Span4Mux_v
    port map (
            O => \N__35921\,
            I => \N__35914\
        );

    \I__7173\ : Span4Mux_v
    port map (
            O => \N__35918\,
            I => \N__35911\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35908\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__35914\,
            I => \N__35904\
        );

    \I__7170\ : Span4Mux_h
    port map (
            O => \N__35911\,
            I => \N__35899\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35899\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35907\,
            I => \N__35896\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__35904\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__35899\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35896\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35889\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__35886\,
            I => \N__35883\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35879\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__35882\,
            I => \N__35876\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__35879\,
            I => \N__35873\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35870\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__35873\,
            I => \N__35865\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35870\,
            I => \N__35865\
        );

    \I__7156\ : Span4Mux_h
    port map (
            O => \N__35865\,
            I => \N__35860\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35857\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35854\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__35860\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35857\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35854\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__7150\ : InMux
    port map (
            O => \N__35847\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__35844\,
            I => \N__35840\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35837\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35834\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35830\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35827\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35824\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__35830\,
            I => \N__35818\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__35827\,
            I => \N__35818\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35824\,
            I => \N__35815\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35812\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__35818\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__35815\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__35812\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35805\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__7135\ : CascadeMux
    port map (
            O => \N__35802\,
            I => \N__35798\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35795\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35792\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__35795\,
            I => \N__35788\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35785\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35782\
        );

    \I__7129\ : Span4Mux_v
    port map (
            O => \N__35788\,
            I => \N__35779\
        );

    \I__7128\ : Span4Mux_h
    port map (
            O => \N__35785\,
            I => \N__35774\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35782\,
            I => \N__35774\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__35779\,
            I => \N__35771\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__35774\,
            I => \N__35768\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__35771\,
            I => \N__35764\
        );

    \I__7123\ : Span4Mux_h
    port map (
            O => \N__35768\,
            I => \N__35761\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35758\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__35764\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__35761\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__35758\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35751\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__7117\ : CascadeMux
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__7116\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35741\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35738\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35734\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35731\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35728\
        );

    \I__7111\ : Span4Mux_v
    port map (
            O => \N__35734\,
            I => \N__35725\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__35731\,
            I => \N__35722\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__35728\,
            I => \N__35719\
        );

    \I__7108\ : Sp12to4
    port map (
            O => \N__35725\,
            I => \N__35715\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__35722\,
            I => \N__35712\
        );

    \I__7106\ : Span4Mux_v
    port map (
            O => \N__35719\,
            I => \N__35709\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35706\
        );

    \I__7104\ : Odrv12
    port map (
            O => \N__35715\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__35712\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__35709\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35706\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35697\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35694\,
            I => \N__35691\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__35691\,
            I => \N__35687\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35684\
        );

    \I__7096\ : Span4Mux_v
    port map (
            O => \N__35687\,
            I => \N__35678\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35678\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35674\
        );

    \I__7093\ : Span4Mux_h
    port map (
            O => \N__35678\,
            I => \N__35671\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35677\,
            I => \N__35668\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35674\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__35671\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__35668\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35661\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__35658\,
            I => \N__35655\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35651\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__35654\,
            I => \N__35648\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35645\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35648\,
            I => \N__35642\
        );

    \I__7082\ : Span4Mux_v
    port map (
            O => \N__35645\,
            I => \N__35636\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35636\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35633\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__35636\,
            I => \N__35629\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35626\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35623\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__35629\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__7075\ : Odrv4
    port map (
            O => \N__35626\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__35623\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35616\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__35613\,
            I => \N__35609\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35606\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35603\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35606\,
            I => \N__35597\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__35603\,
            I => \N__35597\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35594\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__35597\,
            I => \N__35589\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35594\,
            I => \N__35589\
        );

    \I__7064\ : Span4Mux_h
    port map (
            O => \N__35589\,
            I => \N__35585\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35582\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__35585\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35582\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35577\,
            I => \bfn_14_17_0_\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35568\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35568\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35564\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35561\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__35564\,
            I => \N__35556\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35556\
        );

    \I__7053\ : Span4Mux_h
    port map (
            O => \N__35556\,
            I => \N__35552\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35549\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__35552\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__35549\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35544\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35541\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__7047\ : CascadeMux
    port map (
            O => \N__35538\,
            I => \N__35535\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35531\
        );

    \I__7045\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35528\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35524\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__35528\,
            I => \N__35521\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35518\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__35524\,
            I => \N__35515\
        );

    \I__7040\ : Span4Mux_v
    port map (
            O => \N__35521\,
            I => \N__35512\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__35518\,
            I => \N__35509\
        );

    \I__7038\ : Span4Mux_h
    port map (
            O => \N__35515\,
            I => \N__35505\
        );

    \I__7037\ : Span4Mux_h
    port map (
            O => \N__35512\,
            I => \N__35500\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__35509\,
            I => \N__35500\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35497\
        );

    \I__7034\ : Odrv4
    port map (
            O => \N__35505\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__7033\ : Odrv4
    port map (
            O => \N__35500\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35497\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35490\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__7030\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35484\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35484\,
            I => \N__35479\
        );

    \I__7028\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35476\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35473\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35468\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35468\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35465\
        );

    \I__7023\ : Span4Mux_h
    port map (
            O => \N__35468\,
            I => \N__35461\
        );

    \I__7022\ : Span4Mux_v
    port map (
            O => \N__35465\,
            I => \N__35458\
        );

    \I__7021\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35455\
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__35461\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__35458\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35455\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__7017\ : InMux
    port map (
            O => \N__35448\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35445\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__7015\ : InMux
    port map (
            O => \N__35442\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__7014\ : CascadeMux
    port map (
            O => \N__35439\,
            I => \N__35435\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35432\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35428\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35425\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35422\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__35428\,
            I => \N__35417\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__35425\,
            I => \N__35417\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__35422\,
            I => \N__35414\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__35417\,
            I => \N__35408\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__35414\,
            I => \N__35408\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35405\
        );

    \I__7003\ : Odrv4
    port map (
            O => \N__35408\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__35405\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35400\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35397\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35390\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35387\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35383\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35380\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35377\
        );

    \I__6994\ : Span12Mux_v
    port map (
            O => \N__35383\,
            I => \N__35371\
        );

    \I__6993\ : Span12Mux_v
    port map (
            O => \N__35380\,
            I => \N__35371\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35368\
        );

    \I__6991\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35365\
        );

    \I__6990\ : Odrv12
    port map (
            O => \N__35371\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__35368\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__35365\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35358\,
            I => \bfn_14_16_0_\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__35355\,
            I => \N__35352\
        );

    \I__6985\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35348\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35345\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__35348\,
            I => \N__35341\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35338\
        );

    \I__6981\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35335\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__35341\,
            I => \N__35328\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__35338\,
            I => \N__35328\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35335\,
            I => \N__35328\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__35328\,
            I => \N__35324\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35321\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__35324\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__35321\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6973\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35312\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35309\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35306\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__6969\ : Span4Mux_v
    port map (
            O => \N__35306\,
            I => \N__35300\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__35303\,
            I => \N__35297\
        );

    \I__6967\ : Span4Mux_h
    port map (
            O => \N__35300\,
            I => \N__35292\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__35297\,
            I => \N__35289\
        );

    \I__6965\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35284\
        );

    \I__6964\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35284\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__35292\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__35289\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__35284\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35277\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35270\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35267\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35264\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35261\
        );

    \I__6955\ : Span4Mux_v
    port map (
            O => \N__35264\,
            I => \N__35256\
        );

    \I__6954\ : Span4Mux_h
    port map (
            O => \N__35261\,
            I => \N__35253\
        );

    \I__6953\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35248\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35248\
        );

    \I__6951\ : Odrv4
    port map (
            O => \N__35256\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__35253\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__35248\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35241\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35234\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35231\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35228\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__6943\ : Span4Mux_v
    port map (
            O => \N__35228\,
            I => \N__35219\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35219\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35224\,
            I => \N__35216\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__35219\,
            I => \N__35211\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35216\,
            I => \N__35211\
        );

    \I__6938\ : Span4Mux_h
    port map (
            O => \N__35211\,
            I => \N__35207\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35204\
        );

    \I__6936\ : Odrv4
    port map (
            O => \N__35207\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35204\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35199\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__35196\,
            I => \N__35192\
        );

    \I__6932\ : CascadeMux
    port map (
            O => \N__35195\,
            I => \N__35189\
        );

    \I__6931\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35183\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__35183\,
            I => \N__35176\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35173\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__35179\,
            I => \N__35170\
        );

    \I__6925\ : Span4Mux_v
    port map (
            O => \N__35176\,
            I => \N__35165\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35165\
        );

    \I__6923\ : Span4Mux_h
    port map (
            O => \N__35170\,
            I => \N__35161\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__35165\,
            I => \N__35158\
        );

    \I__6921\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35155\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__35161\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__35158\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35155\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6917\ : InMux
    port map (
            O => \N__35148\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35145\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__6915\ : CascadeMux
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__6914\ : InMux
    port map (
            O => \N__35139\,
            I => \N__35135\
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__35138\,
            I => \N__35132\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__35135\,
            I => \N__35128\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35132\,
            I => \N__35125\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35122\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__35128\,
            I => \N__35119\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35114\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35122\,
            I => \N__35114\
        );

    \I__6906\ : Span4Mux_h
    port map (
            O => \N__35119\,
            I => \N__35110\
        );

    \I__6905\ : Span4Mux_v
    port map (
            O => \N__35114\,
            I => \N__35107\
        );

    \I__6904\ : InMux
    port map (
            O => \N__35113\,
            I => \N__35104\
        );

    \I__6903\ : Odrv4
    port map (
            O => \N__35110\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6902\ : Odrv4
    port map (
            O => \N__35107\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__35104\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6900\ : InMux
    port map (
            O => \N__35097\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__6899\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35090\
        );

    \I__6898\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35087\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35081\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__35087\,
            I => \N__35081\
        );

    \I__6895\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35078\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__35081\,
            I => \N__35073\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__35078\,
            I => \N__35073\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__35073\,
            I => \N__35069\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35066\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__35069\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35066\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35061\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__35058\,
            I => \N__35055\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35052\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35047\
        );

    \I__6884\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35042\
        );

    \I__6883\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35042\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__35047\,
            I => \N__35039\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__35042\,
            I => \N__35036\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__35039\,
            I => \N__35032\
        );

    \I__6879\ : Span12Mux_v
    port map (
            O => \N__35036\,
            I => \N__35029\
        );

    \I__6878\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35026\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__35032\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6876\ : Odrv12
    port map (
            O => \N__35029\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__35026\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6874\ : InMux
    port map (
            O => \N__35019\,
            I => \bfn_14_15_0_\
        );

    \I__6873\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35012\
        );

    \I__6872\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35009\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35012\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__35009\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__6869\ : CEMux
    port map (
            O => \N__35004\,
            I => \N__35001\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34998\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__34998\,
            I => \phase_controller_inst2.stoper_hc.N_266_0\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34991\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34987\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34991\,
            I => \N__34984\
        );

    \I__6863\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34981\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__34987\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__34984\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__34981\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6859\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34969\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34966\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34972\,
            I => \N__34963\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34969\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__34966\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__34963\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6853\ : ClkMux
    port map (
            O => \N__34956\,
            I => \N__34953\
        );

    \I__6852\ : GlobalMux
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__6851\ : gio2CtrlBuf
    port map (
            O => \N__34950\,
            I => delay_hc_input_c_g
        );

    \I__6850\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34944\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__34944\,
            I => \N__34941\
        );

    \I__6848\ : Odrv12
    port map (
            O => \N__34941\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__6847\ : CascadeMux
    port map (
            O => \N__34938\,
            I => \N__34934\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34930\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34927\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34924\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34919\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34919\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__34924\,
            I => \N__34914\
        );

    \I__6840\ : Span4Mux_s3_v
    port map (
            O => \N__34919\,
            I => \N__34914\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__34914\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34908\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34901\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34896\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34896\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34893\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34890\
        );

    \I__6832\ : Span12Mux_v
    port map (
            O => \N__34901\,
            I => \N__34887\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34896\,
            I => \phase_controller_inst2.N_139_1\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__34893\,
            I => \phase_controller_inst2.N_139_1\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34890\,
            I => \phase_controller_inst2.N_139_1\
        );

    \I__6828\ : Odrv12
    port map (
            O => \N__34887\,
            I => \phase_controller_inst2.N_139_1\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34875\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34875\,
            I => \phase_controller_inst2.stoper_hc.N_34\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34869\,
            I => \phase_controller_inst2.stoper_hc.m20_nsZ0Z_1\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34860\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34856\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34853\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34850\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__34860\,
            I => \N__34847\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34844\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34856\,
            I => \N__34839\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34839\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34850\,
            I => \N__34836\
        );

    \I__6814\ : Span4Mux_v
    port map (
            O => \N__34847\,
            I => \N__34831\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__34844\,
            I => \N__34831\
        );

    \I__6812\ : Span4Mux_h
    port map (
            O => \N__34839\,
            I => \N__34826\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__34836\,
            I => \N__34826\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__34831\,
            I => \N__34823\
        );

    \I__6809\ : Span4Mux_h
    port map (
            O => \N__34826\,
            I => \N__34820\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__34823\,
            I => \N__34817\
        );

    \I__6807\ : Odrv4
    port map (
            O => \N__34820\,
            I => il_min_comp2_c
        );

    \I__6806\ : Odrv4
    port map (
            O => \N__34817\,
            I => il_min_comp2_c
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34805\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34800\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__34805\,
            I => \N__34796\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34791\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34791\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__34800\,
            I => \N__34788\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34785\
        );

    \I__6797\ : Span4Mux_h
    port map (
            O => \N__34796\,
            I => \N__34780\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34780\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__34788\,
            I => \phase_controller_inst2.stoper_hc.hc_time_passed\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34785\,
            I => \phase_controller_inst2.stoper_hc.hc_time_passed\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__34780\,
            I => \phase_controller_inst2.stoper_hc.hc_time_passed\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34770\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34770\,
            I => \N__34767\
        );

    \I__6790\ : Odrv12
    port map (
            O => \N__34767\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34764\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34758\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34758\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34755\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34747\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34744\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__34750\,
            I => \N__34741\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34747\,
            I => \N__34737\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34744\,
            I => \N__34734\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34731\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34723\
        );

    \I__6778\ : Span4Mux_h
    port map (
            O => \N__34737\,
            I => \N__34713\
        );

    \I__6777\ : Span4Mux_h
    port map (
            O => \N__34734\,
            I => \N__34692\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34692\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34681\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34681\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34681\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34681\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34681\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34723\,
            I => \N__34678\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34667\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34667\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34720\,
            I => \N__34667\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34667\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34667\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34662\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34662\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__34713\,
            I => \N__34659\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34644\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34644\
        );

    \I__6759\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34644\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34644\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34644\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34644\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34644\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34635\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34635\
        );

    \I__6752\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34635\
        );

    \I__6751\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34635\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34624\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34624\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34624\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34624\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34624\
        );

    \I__6745\ : Span4Mux_h
    port map (
            O => \N__34692\,
            I => \N__34619\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34681\,
            I => \N__34619\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__34678\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__34667\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34662\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__34659\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__34644\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34635\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__34624\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__34619\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34602\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34596\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__34596\,
            I => \N__34593\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__34593\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34590\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__6730\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34584\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34581\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__34575\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34572\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34566\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__34566\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34563\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34557\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__34557\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34554\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34548\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__6716\ : Odrv12
    port map (
            O => \N__34545\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34542\,
            I => \bfn_13_20_0_\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34536\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34533\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34527\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__34524\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34521\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34515\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34512\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__34512\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34509\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__34503\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34500\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34494\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34494\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34491\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34485\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__34485\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34482\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__6694\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34476\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__34476\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34473\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34467\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__34467\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34464\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__34458\,
            I => \N__34455\
        );

    \I__6686\ : Odrv12
    port map (
            O => \N__34455\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34452\,
            I => \bfn_13_19_0_\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34446\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__34446\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34443\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__34440\,
            I => \N__34437\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34434\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34431\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__34431\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34428\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34422\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__34422\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34419\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__6673\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34413\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__34413\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34410\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34404\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34401\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__34398\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__6666\ : InMux
    port map (
            O => \N__34395\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__34389\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34386\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34380\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__6659\ : Odrv4
    port map (
            O => \N__34374\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34371\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34365\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34365\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__6655\ : InMux
    port map (
            O => \N__34362\,
            I => \bfn_13_18_0_\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__34356\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34353\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34347\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__34347\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34344\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__6648\ : CascadeMux
    port map (
            O => \N__34341\,
            I => \N__34321\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34308\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34303\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34303\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34300\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34297\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34290\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34290\
        );

    \I__6640\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34290\
        );

    \I__6639\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34279\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34274\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34274\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34269\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34269\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34262\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34262\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34262\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34249\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34249\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34249\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34249\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34249\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34249\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34235\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34315\,
            I => \N__34235\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34232\
        );

    \I__6622\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34229\
        );

    \I__6621\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34226\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34222\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34219\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__34303\,
            I => \N__34216\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34300\,
            I => \N__34209\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__34297\,
            I => \N__34204\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__34290\,
            I => \N__34204\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34199\
        );

    \I__6613\ : InMux
    port map (
            O => \N__34288\,
            I => \N__34199\
        );

    \I__6612\ : CascadeMux
    port map (
            O => \N__34287\,
            I => \N__34187\
        );

    \I__6611\ : CascadeMux
    port map (
            O => \N__34286\,
            I => \N__34184\
        );

    \I__6610\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34169\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34169\
        );

    \I__6608\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34169\
        );

    \I__6607\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34166\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34279\,
            I => \N__34161\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34161\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34154\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34154\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__34249\,
            I => \N__34154\
        );

    \I__6601\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34145\
        );

    \I__6600\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34145\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34145\
        );

    \I__6598\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34145\
        );

    \I__6597\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34134\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34134\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34134\
        );

    \I__6594\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34134\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34134\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34127\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34124\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__34229\,
            I => \N__34119\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34226\,
            I => \N__34119\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34116\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34222\,
            I => \N__34113\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__34219\,
            I => \N__34108\
        );

    \I__6585\ : Span4Mux_v
    port map (
            O => \N__34216\,
            I => \N__34108\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34099\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34099\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34099\
        );

    \I__6581\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34099\
        );

    \I__6580\ : Span12Mux_h
    port map (
            O => \N__34209\,
            I => \N__34092\
        );

    \I__6579\ : Sp12to4
    port map (
            O => \N__34204\,
            I => \N__34092\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__34199\,
            I => \N__34092\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34087\
        );

    \I__6576\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34087\
        );

    \I__6575\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34076\
        );

    \I__6574\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34076\
        );

    \I__6573\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34076\
        );

    \I__6572\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34076\
        );

    \I__6571\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34076\
        );

    \I__6570\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34059\
        );

    \I__6569\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34059\
        );

    \I__6568\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34059\
        );

    \I__6567\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34059\
        );

    \I__6566\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34059\
        );

    \I__6565\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34059\
        );

    \I__6564\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34059\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34059\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34054\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34054\
        );

    \I__6560\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34049\
        );

    \I__6559\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34049\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34042\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34042\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__34161\,
            I => \N__34042\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__34154\,
            I => \N__34035\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__34145\,
            I => \N__34035\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__34134\,
            I => \N__34035\
        );

    \I__6552\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34026\
        );

    \I__6551\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34026\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34026\
        );

    \I__6549\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34026\
        );

    \I__6548\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__34017\
        );

    \I__6547\ : Span4Mux_v
    port map (
            O => \N__34124\,
            I => \N__34017\
        );

    \I__6546\ : Span4Mux_v
    port map (
            O => \N__34119\,
            I => \N__34017\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__34116\,
            I => \N__34017\
        );

    \I__6544\ : Odrv12
    port map (
            O => \N__34113\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__34108\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__34099\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6541\ : Odrv12
    port map (
            O => \N__34092\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__34087\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__34076\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__34059\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__34054\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__34049\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__34042\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6534\ : Odrv4
    port map (
            O => \N__34035\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34026\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__34017\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__33990\,
            I => \N__33972\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__33989\,
            I => \N__33964\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33954\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33954\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__33986\,
            I => \N__33949\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__33985\,
            I => \N__33942\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__33984\,
            I => \N__33938\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__33983\,
            I => \N__33932\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__33982\,
            I => \N__33928\
        );

    \I__6522\ : CascadeMux
    port map (
            O => \N__33981\,
            I => \N__33924\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__33980\,
            I => \N__33921\
        );

    \I__6520\ : CascadeMux
    port map (
            O => \N__33979\,
            I => \N__33917\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__33978\,
            I => \N__33912\
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__33977\,
            I => \N__33908\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__33976\,
            I => \N__33905\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33902\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33899\
        );

    \I__6514\ : CascadeMux
    port map (
            O => \N__33971\,
            I => \N__33892\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__33970\,
            I => \N__33889\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__33969\,
            I => \N__33884\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__33968\,
            I => \N__33880\
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__33967\,
            I => \N__33876\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33860\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__33963\,
            I => \N__33856\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33846\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33846\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33846\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33846\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33954\,
            I => \N__33843\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33838\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33838\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33835\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33828\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33828\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33828\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33825\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33814\
        );

    \I__6494\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33814\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33814\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33814\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33814\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33805\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33805\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33805\
        );

    \I__6487\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33805\
        );

    \I__6486\ : InMux
    port map (
            O => \N__33927\,
            I => \N__33794\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33794\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33794\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33794\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33794\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__33916\,
            I => \N__33790\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33774\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33774\
        );

    \I__6478\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33774\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33769\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33769\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__33902\,
            I => \N__33766\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33759\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__33898\,
            I => \N__33755\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \N__33751\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__33896\,
            I => \N__33747\
        );

    \I__6470\ : InMux
    port map (
            O => \N__33895\,
            I => \N__33739\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33739\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33889\,
            I => \N__33739\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33888\,
            I => \N__33722\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33722\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33722\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33722\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33722\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33722\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33876\,
            I => \N__33722\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33722\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__33874\,
            I => \N__33719\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__33873\,
            I => \N__33715\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33872\,
            I => \N__33711\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__33871\,
            I => \N__33707\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__33870\,
            I => \N__33703\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__33869\,
            I => \N__33699\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__33868\,
            I => \N__33695\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__33867\,
            I => \N__33691\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__33866\,
            I => \N__33687\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__33865\,
            I => \N__33683\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__33864\,
            I => \N__33679\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__33863\,
            I => \N__33675\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33667\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33662\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33856\,
            I => \N__33662\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__33855\,
            I => \N__33658\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33655\
        );

    \I__6442\ : Span4Mux_h
    port map (
            O => \N__33843\,
            I => \N__33650\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__33838\,
            I => \N__33650\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33639\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__33828\,
            I => \N__33639\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33639\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33814\,
            I => \N__33639\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33805\,
            I => \N__33639\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33794\,
            I => \N__33636\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33633\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33630\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__33789\,
            I => \N__33623\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__33788\,
            I => \N__33618\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33611\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33611\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33611\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33606\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33606\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33601\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33601\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33594\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33769\,
            I => \N__33594\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__33766\,
            I => \N__33594\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__33765\,
            I => \N__33590\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__33764\,
            I => \N__33586\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__33763\,
            I => \N__33582\
        );

    \I__6417\ : CascadeMux
    port map (
            O => \N__33762\,
            I => \N__33578\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__33759\,
            I => \N__33575\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33560\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33560\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33560\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33560\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33560\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33560\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33560\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__33739\,
            I => \N__33555\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__33722\,
            I => \N__33555\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33538\
        );

    \I__6405\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33538\
        );

    \I__6404\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33538\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33538\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33538\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33710\,
            I => \N__33538\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33538\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33538\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33521\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33521\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33521\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33521\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33521\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33521\
        );

    \I__6392\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33521\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33521\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33504\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33504\
        );

    \I__6388\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33504\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33504\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33504\
        );

    \I__6385\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33504\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33504\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33504\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__33673\,
            I => \N__33499\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__33672\,
            I => \N__33495\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__33671\,
            I => \N__33491\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33670\,
            I => \N__33485\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__33667\,
            I => \N__33479\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33662\,
            I => \N__33479\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33474\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33474\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__33655\,
            I => \N__33461\
        );

    \I__6373\ : Span4Mux_v
    port map (
            O => \N__33650\,
            I => \N__33461\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__33639\,
            I => \N__33461\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__33636\,
            I => \N__33461\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__33633\,
            I => \N__33461\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33461\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33444\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33444\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33444\
        );

    \I__6365\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33444\
        );

    \I__6364\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33444\
        );

    \I__6363\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33444\
        );

    \I__6362\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33444\
        );

    \I__6361\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33444\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__33611\,
            I => \N__33435\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__33606\,
            I => \N__33435\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__33601\,
            I => \N__33435\
        );

    \I__6357\ : Span4Mux_h
    port map (
            O => \N__33594\,
            I => \N__33435\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33418\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33418\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33418\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33418\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33418\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33418\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33418\
        );

    \I__6349\ : InMux
    port map (
            O => \N__33578\,
            I => \N__33418\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__33575\,
            I => \N__33405\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__33560\,
            I => \N__33405\
        );

    \I__6346\ : Span4Mux_v
    port map (
            O => \N__33555\,
            I => \N__33405\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__33538\,
            I => \N__33405\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33405\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__33504\,
            I => \N__33405\
        );

    \I__6342\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33400\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33400\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33387\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33387\
        );

    \I__6338\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33387\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33387\
        );

    \I__6336\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33387\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33387\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33378\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33378\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33378\
        );

    \I__6331\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33378\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__33479\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33474\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__33461\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__33444\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__33435\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__33418\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__33405\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__33400\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33387\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__33378\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__33357\,
            I => \N__33354\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33351\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33347\
        );

    \I__6317\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33344\
        );

    \I__6316\ : Span4Mux_h
    port map (
            O => \N__33347\,
            I => \N__33340\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__33344\,
            I => \N__33337\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33334\
        );

    \I__6313\ : Sp12to4
    port map (
            O => \N__33340\,
            I => \N__33331\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__33337\,
            I => \N__33328\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33334\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__6310\ : Odrv12
    port map (
            O => \N__33331\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__33328\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__33315\,
            I => \N__33312\
        );

    \I__6305\ : Span4Mux_h
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__6304\ : Span4Mux_v
    port map (
            O => \N__33309\,
            I => \N__33306\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__33306\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33300\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__33294\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__33288\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33281\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33278\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__33281\,
            I => \N__33273\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33273\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__33273\,
            I => \N__33270\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__33270\,
            I => \N__33266\
        );

    \I__6290\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__33266\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33263\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33255\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33252\
        );

    \I__6285\ : Span4Mux_h
    port map (
            O => \N__33252\,
            I => \N__33249\
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__33249\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33243\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__33243\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33237\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__33237\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__33234\,
            I => \N__33229\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33226\
        );

    \I__6277\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33223\
        );

    \I__6276\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33220\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__33226\,
            I => \current_shift_inst.N_1275_i\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__33223\,
            I => \current_shift_inst.N_1275_i\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33220\,
            I => \current_shift_inst.N_1275_i\
        );

    \I__6272\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33210\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33207\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__6269\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33201\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33198\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__33192\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__33186\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__33183\,
            I => \N__33180\
        );

    \I__6261\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33177\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__33177\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33171\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33171\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33168\,
            I => \N__33165\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__33165\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33159\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__33159\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33153\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__33153\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33147\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__33147\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__33141\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33134\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33131\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__33134\,
            I => \N__33127\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33124\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33121\
        );

    \I__6242\ : Odrv12
    port map (
            O => \N__33127\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__33124\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__33121\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33108\,
            I => \N__33105\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__33102\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33099\,
            I => \N__33096\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33096\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__6232\ : InMux
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__33090\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__6230\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33080\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33077\
        );

    \I__6227\ : Span12Mux_h
    port map (
            O => \N__33080\,
            I => \N__33073\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__33077\,
            I => \N__33070\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__33073\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__33070\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33067\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__33060\,
            I => \N__33057\
        );

    \I__6220\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33054\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__6218\ : Span4Mux_v
    port map (
            O => \N__33051\,
            I => \N__33048\
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__33048\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__6216\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33042\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__33042\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33036\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__6212\ : CascadeMux
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__6211\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33027\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__33027\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__33021\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33014\
        );

    \I__6206\ : InMux
    port map (
            O => \N__33017\,
            I => \N__33011\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__33006\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__33006\
        );

    \I__6203\ : Span4Mux_h
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__6202\ : Span4Mux_v
    port map (
            O => \N__33003\,
            I => \N__32998\
        );

    \I__6201\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32993\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32993\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__32998\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32993\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__32982\,
            I => \N__32978\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32975\
        );

    \I__6193\ : Span4Mux_v
    port map (
            O => \N__32978\,
            I => \N__32972\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32969\
        );

    \I__6191\ : Span4Mux_h
    port map (
            O => \N__32972\,
            I => \N__32965\
        );

    \I__6190\ : Span4Mux_h
    port map (
            O => \N__32969\,
            I => \N__32962\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32959\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__32965\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__32962\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32959\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__32952\,
            I => \N__32949\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__6182\ : Span4Mux_v
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__6181\ : Odrv4
    port map (
            O => \N__32940\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__6180\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32934\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__6176\ : Span4Mux_h
    port map (
            O => \N__32925\,
            I => \N__32921\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32918\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__32921\,
            I => \N__32914\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32918\,
            I => \N__32911\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32908\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__32914\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32911\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__32908\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__32898\,
            I => \N__32895\
        );

    \I__6166\ : Span4Mux_h
    port map (
            O => \N__32895\,
            I => \N__32892\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__32892\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32886\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32886\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32877\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32877\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32871\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32868\
        );

    \I__6157\ : Span12Mux_v
    port map (
            O => \N__32868\,
            I => \N__32865\
        );

    \I__6156\ : Odrv12
    port map (
            O => \N__32865\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32859\,
            I => \N__32856\
        );

    \I__6153\ : Span4Mux_v
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__32853\,
            I => \N__32850\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__32850\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32844\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32844\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32838\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__32838\,
            I => \N__32834\
        );

    \I__6146\ : InMux
    port map (
            O => \N__32837\,
            I => \N__32831\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__32834\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32831\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__32826\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32816\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32816\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32813\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32809\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32806\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32803\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__32809\,
            I => \N__32800\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__32806\,
            I => \N__32795\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32795\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__32800\,
            I => \N__32792\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__32795\,
            I => \N__32789\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__32792\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__32789\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32775\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32775\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__32775\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32769\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32764\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32761\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32758\
        );

    \I__6121\ : Span4Mux_v
    port map (
            O => \N__32764\,
            I => \N__32753\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32761\,
            I => \N__32753\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32758\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__32753\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32742\
        );

    \I__6116\ : CascadeMux
    port map (
            O => \N__32747\,
            I => \N__32739\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32736\
        );

    \I__6114\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32733\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32730\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32727\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32724\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32733\,
            I => \N__32717\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__32730\,
            I => \N__32717\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32717\
        );

    \I__6107\ : Span4Mux_h
    port map (
            O => \N__32724\,
            I => \N__32714\
        );

    \I__6106\ : Span4Mux_h
    port map (
            O => \N__32717\,
            I => \N__32711\
        );

    \I__6105\ : Odrv4
    port map (
            O => \N__32714\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__32711\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32703\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32700\
        );

    \I__6101\ : Span4Mux_h
    port map (
            O => \N__32700\,
            I => \N__32697\
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__32697\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__32694\,
            I => \N__32645\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32641\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32634\
        );

    \I__6096\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32634\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32627\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32627\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32627\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32613\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32613\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32613\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32613\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32596\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32596\
        );

    \I__6086\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32596\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32589\
        );

    \I__6084\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32589\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32589\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32578\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32578\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32578\
        );

    \I__6079\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32578\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32578\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32571\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32571\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32571\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32566\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32566\
        );

    \I__6072\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32558\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32551\
        );

    \I__6070\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32551\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32551\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32542\
        );

    \I__6067\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32542\
        );

    \I__6066\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32542\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32542\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32539\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32534\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32534\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32521\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32521\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32521\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32521\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32521\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32521\
        );

    \I__6055\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32510\
        );

    \I__6054\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32510\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32510\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32510\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32510\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32507\
        );

    \I__6049\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32504\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32501\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32498\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32495\
        );

    \I__6045\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32478\
        );

    \I__6044\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32478\
        );

    \I__6043\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32478\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32473\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32473\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32470\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32465\
        );

    \I__6038\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32465\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32460\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32460\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32447\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32447\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32447\
        );

    \I__6032\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32447\
        );

    \I__6031\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32447\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32447\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32442\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32442\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__32578\,
            I => \N__32437\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32571\,
            I => \N__32437\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32434\
        );

    \I__6024\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32427\
        );

    \I__6023\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32427\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32422\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32422\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32419\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32416\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__32551\,
            I => \N__32411\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32411\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32400\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32400\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32400\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32400\
        );

    \I__6012\ : Span4Mux_v
    port map (
            O => \N__32507\,
            I => \N__32400\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32391\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__32501\,
            I => \N__32391\
        );

    \I__6009\ : Span4Mux_v
    port map (
            O => \N__32498\,
            I => \N__32391\
        );

    \I__6008\ : Span4Mux_v
    port map (
            O => \N__32495\,
            I => \N__32391\
        );

    \I__6007\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32377\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32377\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32374\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32365\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32365\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32365\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32365\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32359\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32359\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32356\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32353\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32346\
        );

    \I__5995\ : Span4Mux_h
    port map (
            O => \N__32470\,
            I => \N__32346\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32465\,
            I => \N__32346\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__32460\,
            I => \N__32335\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32335\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__32442\,
            I => \N__32335\
        );

    \I__5990\ : Span4Mux_v
    port map (
            O => \N__32437\,
            I => \N__32335\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__32434\,
            I => \N__32335\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32330\
        );

    \I__5987\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32330\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32427\,
            I => \N__32325\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__32422\,
            I => \N__32325\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__32419\,
            I => \N__32314\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__32416\,
            I => \N__32314\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__32411\,
            I => \N__32314\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__32400\,
            I => \N__32314\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__32391\,
            I => \N__32314\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32303\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32303\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32303\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32303\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32303\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32294\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32294\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32294\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32294\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__32377\,
            I => \N__32287\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32287\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__32365\,
            I => \N__32287\
        );

    \I__5967\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32284\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32359\,
            I => \N__32277\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32277\
        );

    \I__5964\ : Span12Mux_h
    port map (
            O => \N__32353\,
            I => \N__32277\
        );

    \I__5963\ : Span4Mux_h
    port map (
            O => \N__32346\,
            I => \N__32272\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__32335\,
            I => \N__32272\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__32330\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5960\ : Odrv12
    port map (
            O => \N__32325\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__32314\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32303\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__32294\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__32287\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__32284\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5954\ : Odrv12
    port map (
            O => \N__32277\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__32272\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32249\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32245\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32242\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32239\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32245\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5947\ : Odrv12
    port map (
            O => \N__32242\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__32239\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5945\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32227\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32224\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32220\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32227\,
            I => \N__32217\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32214\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32211\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__32220\,
            I => \N__32208\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__32217\,
            I => \N__32205\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__32214\,
            I => \N__32200\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32200\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__32208\,
            I => \N__32195\
        );

    \I__5934\ : Span4Mux_v
    port map (
            O => \N__32205\,
            I => \N__32195\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__32200\,
            I => \N__32192\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__32195\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__32192\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5930\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32181\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32181\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__32181\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__5927\ : CEMux
    port map (
            O => \N__32178\,
            I => \N__32173\
        );

    \I__5926\ : CEMux
    port map (
            O => \N__32177\,
            I => \N__32166\
        );

    \I__5925\ : CEMux
    port map (
            O => \N__32176\,
            I => \N__32163\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32160\
        );

    \I__5923\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32157\
        );

    \I__5922\ : CEMux
    port map (
            O => \N__32171\,
            I => \N__32154\
        );

    \I__5921\ : CEMux
    port map (
            O => \N__32170\,
            I => \N__32151\
        );

    \I__5920\ : CEMux
    port map (
            O => \N__32169\,
            I => \N__32136\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__32166\,
            I => \N__32122\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32122\
        );

    \I__5917\ : Span4Mux_v
    port map (
            O => \N__32160\,
            I => \N__32122\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__32122\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32122\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__32151\,
            I => \N__32119\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32097\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32097\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32097\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32088\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32088\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32088\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32088\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32075\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32075\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32075\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32075\
        );

    \I__5902\ : CEMux
    port map (
            O => \N__32139\,
            I => \N__32071\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32068\
        );

    \I__5900\ : CEMux
    port map (
            O => \N__32135\,
            I => \N__32065\
        );

    \I__5899\ : CEMux
    port map (
            O => \N__32134\,
            I => \N__32062\
        );

    \I__5898\ : CEMux
    port map (
            O => \N__32133\,
            I => \N__32059\
        );

    \I__5897\ : Span4Mux_v
    port map (
            O => \N__32122\,
            I => \N__32056\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__32119\,
            I => \N__32053\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32044\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32044\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32044\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32044\
        );

    \I__5891\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32035\
        );

    \I__5890\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32035\
        );

    \I__5889\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32035\
        );

    \I__5888\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32035\
        );

    \I__5887\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32028\
        );

    \I__5886\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32028\
        );

    \I__5885\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32028\
        );

    \I__5884\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32019\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32019\
        );

    \I__5882\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32019\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32019\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32016\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__32088\,
            I => \N__32013\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32004\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32004\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32004\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32004\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__32075\,
            I => \N__32001\
        );

    \I__5873\ : CEMux
    port map (
            O => \N__32074\,
            I => \N__31998\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__32071\,
            I => \N__31995\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__32068\,
            I => \N__31992\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__32065\,
            I => \N__31981\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__32062\,
            I => \N__31981\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__31981\
        );

    \I__5867\ : Span4Mux_v
    port map (
            O => \N__32056\,
            I => \N__31981\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__32053\,
            I => \N__31981\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__31970\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__31970\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__31970\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__32019\,
            I => \N__31970\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__32016\,
            I => \N__31970\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__32013\,
            I => \N__31963\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31963\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__32001\,
            I => \N__31963\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31960\
        );

    \I__5856\ : Span4Mux_v
    port map (
            O => \N__31995\,
            I => \N__31957\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__31992\,
            I => \N__31954\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__31981\,
            I => \N__31951\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__31970\,
            I => \N__31946\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__31963\,
            I => \N__31946\
        );

    \I__5851\ : Odrv12
    port map (
            O => \N__31960\,
            I => \phase_controller_inst1.m3\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__31957\,
            I => \phase_controller_inst1.m3\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__31954\,
            I => \phase_controller_inst1.m3\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__31951\,
            I => \phase_controller_inst1.m3\
        );

    \I__5847\ : Odrv4
    port map (
            O => \N__31946\,
            I => \phase_controller_inst1.m3\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31932\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__5844\ : Span4Mux_v
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__31926\,
            I => \N__31923\
        );

    \I__5842\ : Span4Mux_h
    port map (
            O => \N__31923\,
            I => \N__31920\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__31920\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31911\,
            I => \N__31906\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31903\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31900\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__31906\,
            I => \N__31897\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31903\,
            I => \N__31894\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31891\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__31897\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5831\ : Odrv12
    port map (
            O => \N__31894\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5830\ : Odrv4
    port map (
            O => \N__31891\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31875\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__31872\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31866\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31862\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__31865\,
            I => \N__31858\
        );

    \I__5821\ : Span12Mux_h
    port map (
            O => \N__31862\,
            I => \N__31855\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31852\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31849\
        );

    \I__5818\ : Odrv12
    port map (
            O => \N__31855\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31852\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31849\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__31842\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31835\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__31838\,
            I => \N__31832\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31829\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31832\,
            I => \N__31826\
        );

    \I__5810\ : Span4Mux_h
    port map (
            O => \N__31829\,
            I => \N__31821\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31826\,
            I => \N__31821\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__31821\,
            I => \N__31818\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__31818\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31812\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31812\,
            I => \N__31807\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31811\,
            I => \N__31802\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31802\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__31807\,
            I => \N__31796\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31793\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__31796\,
            I => \N__31790\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31793\,
            I => \N__31787\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__31790\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__5796\ : Odrv12
    port map (
            O => \N__31787\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31775\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31772\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__31775\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__31772\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31763\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31759\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31763\,
            I => \N__31756\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31753\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31759\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__31756\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31753\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31742\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__31745\,
            I => \N__31737\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__31742\,
            I => \N__31734\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31731\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31728\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31725\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__31734\,
            I => \N__31720\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31720\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31715\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31715\
        );

    \I__5773\ : Span4Mux_h
    port map (
            O => \N__31720\,
            I => \N__31712\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__31715\,
            I => \N__31709\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__31712\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__31709\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__5769\ : CEMux
    port map (
            O => \N__31704\,
            I => \N__31668\
        );

    \I__5768\ : CEMux
    port map (
            O => \N__31703\,
            I => \N__31668\
        );

    \I__5767\ : CEMux
    port map (
            O => \N__31702\,
            I => \N__31668\
        );

    \I__5766\ : CEMux
    port map (
            O => \N__31701\,
            I => \N__31668\
        );

    \I__5765\ : CEMux
    port map (
            O => \N__31700\,
            I => \N__31668\
        );

    \I__5764\ : CEMux
    port map (
            O => \N__31699\,
            I => \N__31668\
        );

    \I__5763\ : CEMux
    port map (
            O => \N__31698\,
            I => \N__31668\
        );

    \I__5762\ : CEMux
    port map (
            O => \N__31697\,
            I => \N__31668\
        );

    \I__5761\ : CEMux
    port map (
            O => \N__31696\,
            I => \N__31668\
        );

    \I__5760\ : CEMux
    port map (
            O => \N__31695\,
            I => \N__31668\
        );

    \I__5759\ : CEMux
    port map (
            O => \N__31694\,
            I => \N__31668\
        );

    \I__5758\ : CEMux
    port map (
            O => \N__31693\,
            I => \N__31668\
        );

    \I__5757\ : GlobalMux
    port map (
            O => \N__31668\,
            I => \N__31665\
        );

    \I__5756\ : gio2CtrlBuf
    port map (
            O => \N__31665\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31656\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31656\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31653\
        );

    \I__5752\ : Odrv12
    port map (
            O => \N__31653\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31641\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31641\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31641\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__31635\,
            I => \N__31632\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__31632\,
            I => \N__31629\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__31629\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31620\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31620\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31620\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__31617\,
            I => \N__31612\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31609\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31604\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31604\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31609\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31604\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__31599\,
            I => \N__31595\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31591\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31588\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31585\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31591\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__31588\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__31585\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31574\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31571\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31574\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31571\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__31566\,
            I => \N__31563\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__31557\,
            I => \N__31554\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__31554\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__31551\,
            I => \N__31548\
        );

    \I__5717\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__31539\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31530\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31530\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31526\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31523\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__31526\,
            I => \N__31520\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__31523\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__31520\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__5705\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31506\
        );

    \I__5704\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31506\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__31506\,
            I => \N__31502\
        );

    \I__5702\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31499\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__31502\,
            I => \N__31496\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__31499\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__31496\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31488\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__31485\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__5695\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__31479\,
            I => \N__31476\
        );

    \I__5693\ : Span4Mux_v
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__5692\ : Span4Mux_h
    port map (
            O => \N__31473\,
            I => \N__31466\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31463\
        );

    \I__5690\ : InMux
    port map (
            O => \N__31471\,
            I => \N__31460\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31455\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31455\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__31466\,
            I => \N__31448\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31448\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__31460\,
            I => \N__31448\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31455\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__31448\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31440\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31436\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31433\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__31436\,
            I => \phase_controller_inst2.un4_running_cry_30_THRU_CO\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31433\,
            I => \phase_controller_inst2.un4_running_cry_30_THRU_CO\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31422\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__31422\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__31419\,
            I => \N__31415\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31410\
        );

    \I__5672\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31410\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__31410\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31398\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31393\
        );

    \I__5667\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31393\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31390\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__31398\,
            I => \N__31387\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__31393\,
            I => \N__31384\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__31390\,
            I => \N__31381\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__31387\,
            I => \N__31378\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__31384\,
            I => \N__31375\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__31381\,
            I => \N__31372\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__31378\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__31375\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__31372\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31359\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__31359\,
            I => \N__31355\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31352\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__31355\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__31352\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31341\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31341\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__5647\ : Span4Mux_h
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__31335\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__31332\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__5644\ : InMux
    port map (
            O => \N__31329\,
            I => \N__31326\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31326\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__31320\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__31314\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31307\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31304\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31307\,
            I => \N__31299\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31299\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__31299\,
            I => \N__31296\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__5632\ : Span4Mux_v
    port map (
            O => \N__31293\,
            I => \N__31290\
        );

    \I__5631\ : Span4Mux_v
    port map (
            O => \N__31290\,
            I => \N__31285\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31282\
        );

    \I__5629\ : InMux
    port map (
            O => \N__31288\,
            I => \N__31279\
        );

    \I__5628\ : Span4Mux_v
    port map (
            O => \N__31285\,
            I => \N__31276\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31282\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__31279\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__31276\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5624\ : ClkMux
    port map (
            O => \N__31269\,
            I => \N__31263\
        );

    \I__5623\ : ClkMux
    port map (
            O => \N__31268\,
            I => \N__31263\
        );

    \I__5622\ : GlobalMux
    port map (
            O => \N__31263\,
            I => \N__31260\
        );

    \I__5621\ : gio2CtrlBuf
    port map (
            O => \N__31260\,
            I => delay_tr_input_c_g
        );

    \I__5620\ : IoInMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5618\ : IoSpan4Mux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5617\ : Span4Mux_s1_v
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__31245\,
            I => s3_phy_c
        );

    \I__5615\ : IoInMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5613\ : Span4Mux_s0_v
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__31233\,
            I => \GB_BUFFER_red_c_g_THRU_CO\
        );

    \I__5611\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31227\,
            I => \phase_controller_inst1.stoper_hc.m34_1\
        );

    \I__5609\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31214\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31214\
        );

    \I__5607\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31214\
        );

    \I__5606\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31210\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__31214\,
            I => \N__31207\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__31213\,
            I => \N__31204\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31210\,
            I => \N__31199\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__31207\,
            I => \N__31199\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31196\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31196\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__31193\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__31185\,
            I => \phase_controller_inst2.stoper_hc.m10Z0Z_1\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31179\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31176\
        );

    \I__5593\ : Span4Mux_v
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__31173\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__31164\,
            I => \N__31161\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__31161\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__5587\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__31155\,
            I => \N__31152\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__31149\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__5583\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31140\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__31137\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__5577\ : Span4Mux_h
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__31125\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__5575\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31119\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31119\,
            I => \N__31116\
        );

    \I__5573\ : Odrv12
    port map (
            O => \N__31116\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__31110\,
            I => \N__31105\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31102\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31099\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__31105\,
            I => \N__31096\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31102\,
            I => \N__31093\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31099\,
            I => \N__31090\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__31096\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__31093\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5563\ : Odrv12
    port map (
            O => \N__31090\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5562\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__31077\,
            I => \N__31074\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__31074\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31068\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__5556\ : Odrv4
    port map (
            O => \N__31065\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__5555\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__31059\,
            I => \N__31056\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__31053\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__31050\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__5550\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__31038\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31032\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__31026\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__5542\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__31014\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__5538\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__31005\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__31002\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__5533\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30987\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__30987\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30981\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__30981\,
            I => \N__30978\
        );

    \I__5527\ : Span4Mux_v
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__5526\ : Span4Mux_h
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__30972\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__5524\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__5522\ : Odrv12
    port map (
            O => \N__30963\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__30951\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30945\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__30939\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30930\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__30930\,
            I => \N__30927\
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__30927\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__5509\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30918\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__30918\,
            I => \N__30915\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__30915\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30909\,
            I => \N__30906\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__30906\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30897\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30897\,
            I => \N__30893\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30890\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__30893\,
            I => \N__30884\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30890\,
            I => \N__30884\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30881\
        );

    \I__5495\ : Span4Mux_v
    port map (
            O => \N__30884\,
            I => \N__30878\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30881\,
            I => \N__30875\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__30878\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__5492\ : Odrv12
    port map (
            O => \N__30875\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__30864\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__5488\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__5486\ : Span4Mux_v
    port map (
            O => \N__30855\,
            I => \N__30852\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__30852\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30846\,
            I => \N__30843\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__30843\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30840\,
            I => \N__30837\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30837\,
            I => \N__30834\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__30834\,
            I => \N__30831\
        );

    \I__5478\ : Odrv4
    port map (
            O => \N__30831\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30828\,
            I => \N__30825\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N__30822\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__30822\,
            I => \N__30819\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__30819\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__30810\,
            I => \N__30807\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__30807\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__30798\,
            I => \N__30795\
        );

    \I__5466\ : Odrv4
    port map (
            O => \N__30795\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__30792\,
            I => \N__30789\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30785\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30782\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30785\,
            I => \N__30779\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__30779\,
            I => \N__30773\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__30776\,
            I => \N__30770\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__30773\,
            I => \N__30766\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__30770\,
            I => \N__30763\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30760\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__30766\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__30763\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30760\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__30744\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30738\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__5446\ : Odrv12
    port map (
            O => \N__30735\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__30723\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30717\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__30714\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30708\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__30702\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__30699\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30692\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30689\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30692\,
            I => \N__30686\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30689\,
            I => \N__30683\
        );

    \I__5429\ : Span4Mux_v
    port map (
            O => \N__30686\,
            I => \N__30680\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__30683\,
            I => \N__30677\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__30680\,
            I => \N__30674\
        );

    \I__5426\ : Sp12to4
    port map (
            O => \N__30677\,
            I => \N__30671\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__30674\,
            I => \N__30668\
        );

    \I__5424\ : Span12Mux_h
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__30668\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5422\ : Odrv12
    port map (
            O => \N__30665\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30657\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30657\,
            I => \N__30654\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__30654\,
            I => \N__30651\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__30651\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__5417\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30645\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30642\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__30639\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__5411\ : Odrv12
    port map (
            O => \N__30630\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__5410\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__5408\ : Span4Mux_h
    port map (
            O => \N__30621\,
            I => \N__30618\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__30618\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30615\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30609\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__30606\,
            I => \N__30602\
        );

    \I__5402\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30599\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__30602\,
            I => \N__30593\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30593\
        );

    \I__5399\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30590\
        );

    \I__5398\ : Sp12to4
    port map (
            O => \N__30593\,
            I => \N__30585\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__30590\,
            I => \N__30585\
        );

    \I__5396\ : Odrv12
    port map (
            O => \N__30585\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30578\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30575\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__30578\,
            I => \N__30572\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30569\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__30572\,
            I => \N__30565\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__30569\,
            I => \N__30562\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30559\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__30565\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__30562\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30559\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30546\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__30543\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30533\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__30536\,
            I => \N__30530\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30533\,
            I => \N__30527\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30524\
        );

    \I__5376\ : Span4Mux_v
    port map (
            O => \N__30527\,
            I => \N__30520\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30517\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30514\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__30520\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5372\ : Odrv12
    port map (
            O => \N__30517\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30514\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__30501\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__30489\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5361\ : Odrv12
    port map (
            O => \N__30480\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__5360\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__5358\ : Odrv12
    port map (
            O => \N__30471\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__5357\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30465\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__30465\,
            I => \N__30462\
        );

    \I__5355\ : Span12Mux_v
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__5354\ : Odrv12
    port map (
            O => \N__30459\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5351\ : Span4Mux_h
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5350\ : Odrv4
    port map (
            O => \N__30447\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__30438\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__30432\,
            I => \N__30429\
        );

    \I__5344\ : Span4Mux_h
    port map (
            O => \N__30429\,
            I => \N__30426\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__30426\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30420\,
            I => \N__30417\
        );

    \I__5340\ : Odrv12
    port map (
            O => \N__30417\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__5337\ : Span4Mux_h
    port map (
            O => \N__30408\,
            I => \N__30403\
        );

    \I__5336\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30400\
        );

    \I__5335\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30397\
        );

    \I__5334\ : Span4Mux_v
    port map (
            O => \N__30403\,
            I => \N__30394\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30391\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30388\
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__30394\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5330\ : Odrv12
    port map (
            O => \N__30391\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__30388\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30375\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__5325\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30368\
        );

    \I__5324\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30365\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30361\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30358\
        );

    \I__5321\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30355\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__30361\,
            I => \N__30352\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__30358\,
            I => \N__30347\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30347\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__30352\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__30347\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__30342\,
            I => \N__30339\
        );

    \I__5314\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__30336\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30333\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30330\,
            I => \N__30326\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30323\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30317\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30317\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30314\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__30317\,
            I => \N__30309\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30309\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__30306\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5302\ : InMux
    port map (
            O => \N__30303\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30300\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30297\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30294\,
            I => \bfn_12_16_0_\
        );

    \I__5298\ : InMux
    port map (
            O => \N__30291\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__30288\,
            I => \N__30284\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30280\
        );

    \I__5295\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30275\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30275\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30280\,
            I => \N__30272\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30267\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__30272\,
            I => \N__30267\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__30264\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__5288\ : InMux
    port map (
            O => \N__30261\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__5287\ : InMux
    port map (
            O => \N__30258\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__5286\ : InMux
    port map (
            O => \N__30255\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30252\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30244\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30241\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30238\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30244\,
            I => \N__30233\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30241\,
            I => \N__30233\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__30238\,
            I => \N__30230\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__30233\,
            I => \N__30227\
        );

    \I__5277\ : Odrv4
    port map (
            O => \N__30230\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__30227\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30222\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30214\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30211\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30208\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30214\,
            I => \N__30205\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__30211\,
            I => \N__30200\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30208\,
            I => \N__30200\
        );

    \I__5268\ : Span12Mux_h
    port map (
            O => \N__30205\,
            I => \N__30197\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__30200\,
            I => \N__30194\
        );

    \I__5266\ : Odrv12
    port map (
            O => \N__30197\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__30194\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30189\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__5263\ : InMux
    port map (
            O => \N__30186\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30183\,
            I => \N__30178\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30175\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30172\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30167\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__30175\,
            I => \N__30167\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30164\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__30167\,
            I => \N__30159\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__30164\,
            I => \N__30159\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__30159\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5253\ : InMux
    port map (
            O => \N__30156\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30153\,
            I => \bfn_12_15_0_\
        );

    \I__5251\ : InMux
    port map (
            O => \N__30150\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__5250\ : InMux
    port map (
            O => \N__30147\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__5249\ : InMux
    port map (
            O => \N__30144\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30141\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__30138\,
            I => \N__30135\
        );

    \I__5246\ : InMux
    port map (
            O => \N__30135\,
            I => \N__30130\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30127\
        );

    \I__5244\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30124\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30121\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30116\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30124\,
            I => \N__30116\
        );

    \I__5240\ : Span4Mux_v
    port map (
            O => \N__30121\,
            I => \N__30113\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__30116\,
            I => \N__30110\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__30113\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__30110\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30105\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30097\
        );

    \I__5234\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30094\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30091\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__30097\,
            I => \N__30088\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30083\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30083\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__30088\,
            I => \N__30080\
        );

    \I__5228\ : Span4Mux_v
    port map (
            O => \N__30083\,
            I => \N__30077\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__30080\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__30077\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5225\ : InMux
    port map (
            O => \N__30072\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30069\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30061\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30058\
        );

    \I__5221\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30055\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30061\,
            I => \N__30052\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__30049\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__30055\,
            I => \N__30044\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__30052\,
            I => \N__30044\
        );

    \I__5216\ : Span4Mux_h
    port map (
            O => \N__30049\,
            I => \N__30041\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__30044\,
            I => \N__30038\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__30041\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__30038\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5212\ : InMux
    port map (
            O => \N__30033\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__5211\ : InMux
    port map (
            O => \N__30030\,
            I => \bfn_12_14_0_\
        );

    \I__5210\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30020\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__30023\,
            I => \N__30017\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__30020\,
            I => \N__30013\
        );

    \I__5206\ : InMux
    port map (
            O => \N__30017\,
            I => \N__30008\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30016\,
            I => \N__30008\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__30013\,
            I => \N__30005\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__30008\,
            I => \N__30002\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__30005\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__30002\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5200\ : InMux
    port map (
            O => \N__29997\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29994\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29971\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29971\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29971\
        );

    \I__5195\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29971\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29962\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29962\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29962\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29962\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29934\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29934\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29934\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29934\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29971\,
            I => \N__29929\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29929\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29922\
        );

    \I__5183\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29922\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29922\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29913\
        );

    \I__5180\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29913\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29913\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29913\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29909\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29900\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29900\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29900\
        );

    \I__5173\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29900\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29893\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29893\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29893\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29884\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29884\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29884\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29884\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29881\
        );

    \I__5164\ : Sp12to4
    port map (
            O => \N__29929\,
            I => \N__29874\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29874\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29913\,
            I => \N__29874\
        );

    \I__5161\ : IoInMux
    port map (
            O => \N__29912\,
            I => \N__29871\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29909\,
            I => \N__29858\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29858\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29893\,
            I => \N__29858\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29884\,
            I => \N__29858\
        );

    \I__5156\ : Span12Mux_h
    port map (
            O => \N__29881\,
            I => \N__29858\
        );

    \I__5155\ : Span12Mux_v
    port map (
            O => \N__29874\,
            I => \N__29858\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29855\
        );

    \I__5153\ : Odrv12
    port map (
            O => \N__29858\,
            I => \phase_controller_inst2.m3_0\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__29855\,
            I => \phase_controller_inst2.m3_0\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29850\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__29847\,
            I => \N__29843\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29838\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29838\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29834\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29831\
        );

    \I__5145\ : Span4Mux_h
    port map (
            O => \N__29834\,
            I => \N__29828\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29831\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__29828\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29817\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__29817\,
            I => \N__29813\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29810\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__29813\,
            I => \N__29803\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29803\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29800\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29797\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__29803\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__29800\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__29797\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__29790\,
            I => \N__29787\
        );

    \I__5130\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__5127\ : Span4Mux_h
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__29775\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__5125\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29769\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29769\,
            I => \N__29765\
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__29768\,
            I => \N__29762\
        );

    \I__5122\ : Span4Mux_v
    port map (
            O => \N__29765\,
            I => \N__29757\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29750\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29750\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29750\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__29757\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29750\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__5113\ : Span4Mux_v
    port map (
            O => \N__29736\,
            I => \N__29733\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__29733\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29727\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__5109\ : Span12Mux_v
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__5108\ : Odrv12
    port map (
            O => \N__29721\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29715\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29706\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__29703\,
            I => \N__29698\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29693\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29693\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__29698\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29693\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29681\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29677\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29674\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29671\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29677\,
            I => \N__29668\
        );

    \I__5091\ : Span4Mux_v
    port map (
            O => \N__29674\,
            I => \N__29665\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29662\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__29668\,
            I => \N__29657\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__29665\,
            I => \N__29657\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__29662\,
            I => \N__29654\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__29657\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__29654\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29649\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29646\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__29643\,
            I => \N__29639\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29634\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29634\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29631\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__29631\,
            I => \N__29627\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29624\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__29627\,
            I => \N__29621\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__29624\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__29621\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29616\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__29613\,
            I => \N__29609\
        );

    \I__5071\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29605\
        );

    \I__5070\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29602\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29599\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29594\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29602\,
            I => \N__29594\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__29599\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5065\ : Odrv12
    port map (
            O => \N__29594\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29589\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__29586\,
            I => \N__29582\
        );

    \I__5062\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29578\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29575\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29572\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__29578\,
            I => \N__29567\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__29575\,
            I => \N__29567\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29572\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5056\ : Odrv12
    port map (
            O => \N__29567\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5055\ : InMux
    port map (
            O => \N__29562\,
            I => \bfn_12_11_0_\
        );

    \I__5054\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29552\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29552\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29549\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__29552\,
            I => \N__29546\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__29549\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5049\ : Odrv12
    port map (
            O => \N__29546\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29541\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__29538\,
            I => \N__29534\
        );

    \I__5046\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29529\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29529\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29525\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29522\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__29525\,
            I => \N__29519\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__29522\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__29519\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29514\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29504\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29504\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29501\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__29504\,
            I => \N__29498\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__29501\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__29498\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29493\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__29490\,
            I => \N__29486\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29480\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29480\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29477\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__29480\,
            I => \N__29474\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29477\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__29474\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__5024\ : InMux
    port map (
            O => \N__29469\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29459\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29459\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29456\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29453\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29456\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__29453\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29448\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__5016\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29441\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29438\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29435\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29438\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__29435\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29430\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29424\,
            I => \N__29420\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29417\
        );

    \I__5007\ : Span4Mux_h
    port map (
            O => \N__29420\,
            I => \N__29414\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__29417\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__29414\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5004\ : InMux
    port map (
            O => \N__29409\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29406\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__5002\ : InMux
    port map (
            O => \N__29403\,
            I => \bfn_12_10_0_\
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__29400\,
            I => \N__29396\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29391\
        );

    \I__4999\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29391\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29391\,
            I => \N__29387\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29384\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__29387\,
            I => \N__29381\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__29384\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__29381\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29376\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29366\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29366\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29363\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29360\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__29363\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__29360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29355\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__4985\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29346\
        );

    \I__4984\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29346\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29342\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29339\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__29342\,
            I => \N__29336\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__29339\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__29336\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29331\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__29328\,
            I => \N__29324\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29319\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29319\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29315\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29312\
        );

    \I__4972\ : Span4Mux_v
    port map (
            O => \N__29315\,
            I => \N__29309\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__29312\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__29309\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4969\ : InMux
    port map (
            O => \N__29304\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29295\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29295\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29295\,
            I => \N__29291\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29288\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__29291\,
            I => \N__29285\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29288\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__29285\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4961\ : InMux
    port map (
            O => \N__29280\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__4960\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__29274\,
            I => \N__29270\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29267\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__29264\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4954\ : InMux
    port map (
            O => \N__29259\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29249\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__29249\,
            I => \N__29243\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29246\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__29243\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29238\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29228\
        );

    \I__4944\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29225\
        );

    \I__4943\ : Span4Mux_h
    port map (
            O => \N__29228\,
            I => \N__29222\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29225\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__29222\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4940\ : InMux
    port map (
            O => \N__29217\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__4939\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__29207\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__29204\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4934\ : InMux
    port map (
            O => \N__29199\,
            I => \bfn_12_9_0_\
        );

    \I__4933\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29192\
        );

    \I__4932\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__29189\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__29186\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29181\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29174\
        );

    \I__4926\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29171\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29168\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__29171\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__29168\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29163\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29156\
        );

    \I__4920\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29150\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29153\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__29150\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29145\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__4915\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29139\,
            I => \N__29135\
        );

    \I__4913\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29132\
        );

    \I__4912\ : Span4Mux_v
    port map (
            O => \N__29135\,
            I => \N__29129\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29132\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__29129\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4909\ : InMux
    port map (
            O => \N__29124\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__4908\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29117\
        );

    \I__4907\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29109\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29109\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__29109\,
            I => \N__29106\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__29106\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29099\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29096\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__29099\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29096\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4898\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29088\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__29088\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29081\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29078\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29081\,
            I => \N__29075\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__29078\,
            I => \N__29069\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__29075\,
            I => \N__29066\
        );

    \I__4891\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29059\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29059\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29059\
        );

    \I__4888\ : Odrv12
    port map (
            O => \N__29069\,
            I => \phase_controller_inst1.start_latched\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__29066\,
            I => \phase_controller_inst1.start_latched\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__29059\,
            I => \phase_controller_inst1.start_latched\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__29052\,
            I => \N__29049\
        );

    \I__4884\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29043\
        );

    \I__4883\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29043\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__29040\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__4880\ : InMux
    port map (
            O => \N__29037\,
            I => \N__29031\
        );

    \I__4879\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29031\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__4876\ : Span4Mux_h
    port map (
            O => \N__29025\,
            I => \N__29022\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__29022\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__29016\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__4872\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29009\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29005\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__29002\
        );

    \I__4869\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28999\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__29005\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__29002\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28999\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28989\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__28989\,
            I => \N__28985\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__28985\,
            I => \phase_controller_inst2.N_38\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28982\,
            I => \phase_controller_inst2.N_38\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28974\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28970\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28967\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__28970\,
            I => \N__28964\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__28967\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__28964\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28959\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__28956\,
            I => \N__28952\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__28955\,
            I => \N__28949\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28944\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28944\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28944\,
            I => \phase_controller_inst2.stoper_tr.N_38_i\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28937\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28934\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28931\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28934\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__28931\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28926\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28919\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28922\,
            I => \N__28916\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28919\,
            I => \N__28913\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__28916\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__28913\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28908\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__4836\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28901\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28898\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28901\,
            I => \N__28895\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28898\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__28895\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28890\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28881\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__28881\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28874\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28870\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28867\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28864\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28861\
        );

    \I__4822\ : Span12Mux_v
    port map (
            O => \N__28867\,
            I => \N__28858\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28864\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4820\ : Odrv12
    port map (
            O => \N__28861\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4819\ : Odrv12
    port map (
            O => \N__28858\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28848\,
            I => \N__28843\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28840\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28836\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__28843\,
            I => \N__28833\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__28840\,
            I => \N__28830\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28827\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28824\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__28833\,
            I => \N__28817\
        );

    \I__4809\ : Span4Mux_v
    port map (
            O => \N__28830\,
            I => \N__28817\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28817\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__28824\,
            I => \N__28814\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__28817\,
            I => \N__28811\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__28814\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__28811\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28798\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28795\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28792\
        );

    \I__4799\ : Span4Mux_h
    port map (
            O => \N__28798\,
            I => \N__28789\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28786\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__28792\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__28789\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4795\ : Odrv12
    port map (
            O => \N__28786\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28779\,
            I => \N__28775\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28771\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28775\,
            I => \N__28768\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28765\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28761\
        );

    \I__4789\ : Span4Mux_h
    port map (
            O => \N__28768\,
            I => \N__28756\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28765\,
            I => \N__28756\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28753\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__28761\,
            I => \N__28750\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__28756\,
            I => \N__28745\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__28753\,
            I => \N__28745\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__28750\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__28745\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28734\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28734\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__4778\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28728\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__28719\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28710\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28707\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__28704\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28698\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28698\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__4766\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28691\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__28694\,
            I => \N__28688\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28691\,
            I => \N__28685\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28682\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__28685\,
            I => \N__28678\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28675\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28669\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__28678\,
            I => \N__28664\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__28675\,
            I => \N__28664\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28659\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28659\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28656\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28653\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__28664\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28659\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28656\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4750\ : Odrv12
    port map (
            O => \N__28653\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28638\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28635\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__28635\,
            I => \N__28632\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__28632\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__28629\,
            I => \N__28625\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28621\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28616\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28616\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28621\,
            I => \N__28611\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__28616\,
            I => \N__28611\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__28596\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4732\ : IoInMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__4730\ : Span4Mux_s1_v
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__4729\ : Span4Mux_h
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__28581\,
            I => s4_phy_c
        );

    \I__4727\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28575\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__4725\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28569\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28569\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28560\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__4720\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__28554\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28545\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28545\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28539\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28530\,
            I => \N__28527\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__28527\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28521\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28512\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__28512\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__4703\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28503\,
            I => \N__28500\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__28500\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__4700\ : CascadeMux
    port map (
            O => \N__28497\,
            I => \N__28494\
        );

    \I__4699\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28488\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28488\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28484\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28481\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__28484\,
            I => \N__28478\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__28481\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__28478\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28473\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28464\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28464\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__28464\,
            I => \N__28460\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28457\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__28460\,
            I => \N__28454\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__28457\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__28454\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28449\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28440\
        );

    \I__4682\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28440\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28436\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28433\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__28436\,
            I => \N__28430\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28433\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__28430\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28425\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__28419\,
            I => \N__28414\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28411\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28408\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__28414\,
            I => \N__28403\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__28411\,
            I => \N__28403\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__28408\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__28403\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4667\ : InMux
    port map (
            O => \N__28398\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__4666\ : InMux
    port map (
            O => \N__28395\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28388\
        );

    \I__4664\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28385\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28381\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28378\
        );

    \I__4661\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28375\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__28381\,
            I => \N__28372\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__28378\,
            I => \N__28369\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28375\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__28372\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__28369\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28359\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28359\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28356\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28353\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__28350\,
            I => \N__28346\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28341\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28346\,
            I => \N__28341\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28337\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28334\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__28331\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28326\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28317\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28317\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__28317\,
            I => \N__28313\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28310\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__28313\,
            I => \N__28307\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28310\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__28307\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28302\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28290\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28286\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28283\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__28286\,
            I => \N__28280\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__28283\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__28280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28275\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28266\
        );

    \I__4624\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28266\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28262\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__28262\,
            I => \N__28256\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__28259\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__28256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28251\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__28248\,
            I => \N__28244\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__28247\,
            I => \N__28241\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28236\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28236\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28236\,
            I => \N__28232\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28235\,
            I => \N__28229\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__28232\,
            I => \N__28226\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__28229\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__28226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28221\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28218\,
            I => \N__28212\
        );

    \I__4606\ : InMux
    port map (
            O => \N__28217\,
            I => \N__28212\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__28212\,
            I => \N__28208\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28205\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__28208\,
            I => \N__28202\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28205\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__28202\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28197\,
            I => \bfn_11_15_0_\
        );

    \I__4599\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28187\
        );

    \I__4598\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28187\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28184\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__28187\,
            I => \N__28181\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__28184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__28181\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28176\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__4592\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28169\
        );

    \I__4591\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28166\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__28169\,
            I => \N__28163\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28166\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__28163\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4587\ : InMux
    port map (
            O => \N__28158\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__4586\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28151\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28145\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__28148\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4582\ : Odrv12
    port map (
            O => \N__28145\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28140\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__4580\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28133\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28130\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28127\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__28130\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__28127\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28122\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__4574\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28115\
        );

    \I__4573\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28112\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__28115\,
            I => \N__28109\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__28112\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__28109\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4569\ : InMux
    port map (
            O => \N__28104\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__4568\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28097\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28094\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__28097\,
            I => \N__28091\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__28094\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__28091\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4563\ : InMux
    port map (
            O => \N__28086\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__4562\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28079\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28076\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28073\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__28076\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4558\ : Odrv12
    port map (
            O => \N__28073\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4557\ : InMux
    port map (
            O => \N__28068\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \N__28061\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__28064\,
            I => \N__28058\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28053\
        );

    \I__4553\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28053\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28049\
        );

    \I__4551\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28046\
        );

    \I__4550\ : Sp12to4
    port map (
            O => \N__28049\,
            I => \N__28043\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__28046\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__28043\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28038\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28029\
        );

    \I__4545\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28029\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__28029\,
            I => \N__28025\
        );

    \I__4543\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28022\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__28025\,
            I => \N__28019\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__28022\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__28019\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4539\ : InMux
    port map (
            O => \N__28014\,
            I => \bfn_11_14_0_\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28007\
        );

    \I__4537\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28004\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__28001\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__28004\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__28001\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27996\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__27993\,
            I => \N__27989\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__27992\,
            I => \N__27986\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27981\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27981\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27981\,
            I => \phase_controller_inst1.stoper_tr.N_42_i\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27974\
        );

    \I__4526\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27971\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27974\,
            I => \N__27968\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27971\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__27968\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27963\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27956\
        );

    \I__4520\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27953\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27956\,
            I => \N__27950\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__27953\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__27950\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27945\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27938\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27935\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27938\,
            I => \N__27932\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__27935\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__27932\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27927\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27920\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27923\,
            I => \N__27917\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27920\,
            I => \N__27914\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__27917\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__27914\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27909\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27902\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27899\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27896\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__27899\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4499\ : Odrv12
    port map (
            O => \N__27896\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27891\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27888\,
            I => \N__27884\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27881\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27878\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27881\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__27878\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27873\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27866\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27863\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__27866\,
            I => \N__27860\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27863\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__27860\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27855\,
            I => \bfn_11_13_0_\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27849\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__27846\,
            I => \N__27843\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__27843\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__27840\,
            I => \N__27837\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27834\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27831\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__27828\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27822\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__27816\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__27807\,
            I => \N__27804\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__27801\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__4467\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27795\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27795\,
            I => \N__27792\
        );

    \I__4465\ : Odrv12
    port map (
            O => \N__27792\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__27789\,
            I => \N__27786\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27780\
        );

    \I__4461\ : Odrv12
    port map (
            O => \N__27780\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27774\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__27774\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27765\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27759\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27759\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27756\,
            I => \N__27753\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27750\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__27750\,
            I => \N__27747\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__27747\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27741\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27741\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27732\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27732\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27729\,
            I => \phase_controller_inst1.un4_running_cry_30\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27726\,
            I => \N__27720\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27720\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27720\,
            I => \phase_controller_inst1.un4_running_cry_30_THRU_CO\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27714\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27714\,
            I => \N__27711\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__27711\,
            I => \phase_controller_inst1.N_42\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27704\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27700\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27697\
        );

    \I__4434\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27694\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__27700\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__27697\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__27694\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4430\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__27678\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27669\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__27657\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__4418\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__27648\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__27639\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__27636\,
            I => \N__27633\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27630\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27624\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27621\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__27618\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__27615\,
            I => \N__27612\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27609\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27609\,
            I => \N__27606\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__27606\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__27603\,
            I => \N__27600\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27597\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27597\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__4398\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27588\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27585\
        );

    \I__4396\ : Odrv12
    port map (
            O => \N__27585\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27582\,
            I => \N__27579\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27579\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27573\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__27573\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__27570\,
            I => \N__27567\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27564\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27564\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27558\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27555\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__27555\,
            I => \N__27552\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__27552\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__27549\,
            I => \N__27546\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27543\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27543\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27534\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__27534\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__4377\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__27525\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27519\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__27516\,
            I => \N__27513\
        );

    \I__4372\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__27510\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__27498\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27492\,
            I => \N__27489\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27489\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__4363\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__27480\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4359\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__27468\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__4354\ : Odrv12
    port map (
            O => \N__27459\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27450\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27450\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__4350\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27444\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__27441\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27435\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27432\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27426\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__4342\ : Odrv12
    port map (
            O => \N__27423\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__27420\,
            I => \N__27417\
        );

    \I__4340\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27414\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__4338\ : InMux
    port map (
            O => \N__27411\,
            I => \phase_controller_inst2.un4_running_cry_30\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__27405\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27393\
        );

    \I__4333\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27393\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__27393\,
            I => \N__27390\
        );

    \I__4331\ : Odrv12
    port map (
            O => \N__27390\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__27387\,
            I => \N__27384\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__27381\,
            I => \N__27378\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__27378\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27372\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__27369\,
            I => \N__27366\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27360\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27360\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4320\ : Span4Mux_h
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__27354\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__27351\,
            I => \N__27348\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27345\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__4315\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27337\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27334\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27331\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27328\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__27334\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27331\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4309\ : Odrv12
    port map (
            O => \N__27328\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__4308\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27318\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27313\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__27317\,
            I => \N__27309\
        );

    \I__4305\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27306\
        );

    \I__4304\ : Span4Mux_v
    port map (
            O => \N__27313\,
            I => \N__27303\
        );

    \I__4303\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27298\
        );

    \I__4302\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27298\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__27306\,
            I => \N__27295\
        );

    \I__4300\ : Span4Mux_h
    port map (
            O => \N__27303\,
            I => \N__27290\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27290\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__27295\,
            I => \N__27287\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__27290\,
            I => \N__27284\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__27287\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__27284\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__4294\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27273\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27273\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27273\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27267\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__27267\,
            I => \N__27264\
        );

    \I__4289\ : Odrv12
    port map (
            O => \N__27264\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__4287\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__27255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27249\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27237\
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__27237\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27231\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__4276\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__27222\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__27213\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4270\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27204\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4266\ : Span12Mux_h
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__4265\ : Odrv12
    port map (
            O => \N__27192\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__27183\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__4261\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__27171\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__27162\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__4254\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__27156\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__4252\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27147\
        );

    \I__4250\ : Odrv12
    port map (
            O => \N__27147\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__4248\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27138\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__4244\ : Span4Mux_h
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__27126\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__27114\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__4238\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__27102\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27093\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__27093\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27084\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__27084\,
            I => \N__27081\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__27081\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__4226\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27072\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__27072\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27066\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27066\,
            I => \N__27063\
        );

    \I__4222\ : Odrv12
    port map (
            O => \N__27063\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__4220\ : InMux
    port map (
            O => \N__27057\,
            I => \N__27054\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__27054\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__4218\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27048\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27048\,
            I => \N__27045\
        );

    \I__4216\ : Odrv12
    port map (
            O => \N__27045\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__4214\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27036\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__27036\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__4211\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__27024\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__4208\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__27015\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__4205\ : InMux
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__27009\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__27006\,
            I => \N__27003\
        );

    \I__4202\ : InMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27000\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__26994\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__26991\,
            I => \N__26988\
        );

    \I__4197\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26985\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26985\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__26979\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__26976\,
            I => \N__26973\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26970\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26961\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__26961\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__26958\,
            I => \N__26955\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26952\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__26946\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__26937\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__4179\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26931\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26922\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26913\,
            I => \N__26910\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__26907\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26898\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__26889\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__26877\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26868\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26862\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__4152\ : Odrv12
    port map (
            O => \N__26853\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26844\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__26844\,
            I => \N__26841\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__26841\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26835\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__4143\ : Odrv12
    port map (
            O => \N__26826\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__26820\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26814\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26814\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__26805\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__26793\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26787\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__26778\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__26772\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26766\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__26757\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26748\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__26748\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__26739\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__26736\,
            I => \N__26733\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26730\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__26718\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__26709\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__26706\,
            I => \N__26703\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26700\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__26691\,
            I => \N__26688\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__26688\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__26679\,
            I => \N__26676\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__26676\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__26667\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__4087\ : Sp12to4
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__4086\ : Odrv12
    port map (
            O => \N__26655\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__26652\,
            I => \N__26649\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__26637\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__26625\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__4073\ : Span12Mux_v
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__26613\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__4071\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26606\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26601\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26598\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26593\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26593\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26601\,
            I => \N__26590\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__26598\,
            I => \N__26587\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__26593\,
            I => \N__26584\
        );

    \I__4063\ : Span4Mux_v
    port map (
            O => \N__26590\,
            I => \N__26581\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__26587\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4061\ : Odrv12
    port map (
            O => \N__26584\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26581\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__26574\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26565\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26565\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__26565\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26558\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26558\,
            I => \N__26550\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26555\,
            I => \N__26550\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__26550\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__26547\,
            I => \N__26543\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__26546\,
            I => \N__26540\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26537\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26531\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26534\,
            I => \N__26528\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__26531\,
            I => \N__26525\
        );

    \I__4043\ : Span4Mux_v
    port map (
            O => \N__26528\,
            I => \N__26522\
        );

    \I__4042\ : Span4Mux_v
    port map (
            O => \N__26525\,
            I => \N__26519\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__26522\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__26519\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__4036\ : Span4Mux_h
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__26502\,
            I => \N__26499\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__26499\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__26496\,
            I => \N__26493\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26490\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26490\,
            I => \N__26487\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__26487\,
            I => \N__26484\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__26484\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__26481\,
            I => \N__26478\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__26469\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__4022\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26460\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__26460\,
            I => \N__26457\
        );

    \I__4020\ : Span4Mux_v
    port map (
            O => \N__26457\,
            I => \N__26454\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__26454\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__26451\,
            I => \N__26448\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26445\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__26442\,
            I => \N__26439\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__26439\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26433\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__26433\,
            I => \N__26430\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__26430\,
            I => \N__26427\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__26427\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__26424\,
            I => \phase_controller_inst1.N_42_cascade_\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26412\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26412\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__26412\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__26409\,
            I => \N__26405\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__26408\,
            I => \N__26402\
        );

    \I__4002\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26397\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26397\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26397\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26390\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26386\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26383\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26380\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26386\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__26383\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__26380\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26364\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26361\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26358\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26355\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__26364\,
            I => \N__26350\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26350\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26347\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__26355\,
            I => \N__26344\
        );

    \I__3983\ : Span4Mux_v
    port map (
            O => \N__26350\,
            I => \N__26341\
        );

    \I__3982\ : Span4Mux_h
    port map (
            O => \N__26347\,
            I => \N__26336\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__26344\,
            I => \N__26336\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__26341\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3979\ : Odrv4
    port map (
            O => \N__26336\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__26331\,
            I => \N__26328\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26322\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26322\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__26322\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__3974\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26315\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26312\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26315\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26312\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__26307\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__3969\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26298\
        );

    \I__3968\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26298\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__26298\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26289\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26289\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__26289\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26283\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26283\,
            I => \phase_controller_inst1.N_43\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__26280\,
            I => \phase_controller_inst1.N_43_cascade_\
        );

    \I__3960\ : CEMux
    port map (
            O => \N__26277\,
            I => \N__26274\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__26274\,
            I => \N__26271\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__26271\,
            I => \phase_controller_inst1.stoper_tr.N_43_0\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__26268\,
            I => \N__26263\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__26267\,
            I => \N__26260\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26253\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26253\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26253\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26253\,
            I => \phase_controller_inst1.running\
        );

    \I__3951\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26242\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26239\
        );

    \I__3948\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26236\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__26242\,
            I => \N__26233\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26230\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__26236\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__26233\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3943\ : Odrv12
    port map (
            O => \N__26230\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26219\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26216\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26211\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26208\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26203\
        );

    \I__3937\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26203\
        );

    \I__3936\ : Span4Mux_h
    port map (
            O => \N__26211\,
            I => \N__26200\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__26208\,
            I => \N__26197\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26194\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__26200\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__26197\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__26194\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__3930\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26184\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__26184\,
            I => \N__26180\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26177\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__26180\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26177\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26169\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26169\,
            I => \N__26164\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26159\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26159\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__26164\,
            I => \N__26153\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__26159\,
            I => \N__26153\
        );

    \I__3919\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26150\
        );

    \I__3918\ : Span4Mux_h
    port map (
            O => \N__26153\,
            I => \N__26147\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__26150\,
            I => \N__26144\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__26147\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__3915\ : Odrv12
    port map (
            O => \N__26144\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__26139\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__3912\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26127\
        );

    \I__3911\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26127\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26127\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26121\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26117\
        );

    \I__3907\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26114\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__26117\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__26114\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__3904\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26104\
        );

    \I__3903\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26099\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26107\,
            I => \N__26099\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__26104\,
            I => \N__26096\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26092\
        );

    \I__3899\ : Span4Mux_h
    port map (
            O => \N__26096\,
            I => \N__26089\
        );

    \I__3898\ : InMux
    port map (
            O => \N__26095\,
            I => \N__26086\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__26092\,
            I => \N__26083\
        );

    \I__3896\ : Sp12to4
    port map (
            O => \N__26089\,
            I => \N__26078\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26078\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__26083\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__3893\ : Odrv12
    port map (
            O => \N__26078\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__26073\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26064\
        );

    \I__3890\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26064\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__26064\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__26054\
        );

    \I__3886\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26051\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__26054\,
            I => \N__26047\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__26051\,
            I => \N__26044\
        );

    \I__3883\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26041\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__26047\,
            I => \N__26036\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__26044\,
            I => \N__26036\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__26041\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__26036\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__3878\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26028\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__26028\,
            I => \N__26024\
        );

    \I__3876\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26021\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__26024\,
            I => \N__26015\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26015\
        );

    \I__3873\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26012\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__26015\,
            I => \N__26008\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26005\
        );

    \I__3870\ : InMux
    port map (
            O => \N__26011\,
            I => \N__26002\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__26008\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__3868\ : Odrv12
    port map (
            O => \N__26005\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__26002\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25992\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25988\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25984\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__25988\,
            I => \N__25981\
        );

    \I__3862\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25978\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25984\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25981\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__25978\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25967\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25963\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25960\
        );

    \I__3855\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25957\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25953\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__25960\,
            I => \N__25950\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25947\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__25956\,
            I => \N__25944\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__25953\,
            I => \N__25937\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__25950\,
            I => \N__25937\
        );

    \I__3848\ : Span4Mux_v
    port map (
            O => \N__25947\,
            I => \N__25937\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25934\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__25937\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__25934\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25923\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25923\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25923\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__25920\,
            I => \N__25917\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25911\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25911\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25911\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25903\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25900\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25897\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25903\,
            I => \N__25891\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25891\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25897\,
            I => \N__25888\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25885\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__25891\,
            I => \N__25882\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__25888\,
            I => \N__25877\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25885\,
            I => \N__25877\
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__25882\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__25877\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25868\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25864\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25861\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25858\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25864\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__3820\ : Odrv12
    port map (
            O => \N__25861\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25858\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25845\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25845\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25845\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25833\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25833\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__25833\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25830\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25827\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25824\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25821\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25818\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25812\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25812\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__3802\ : Glb2LocalMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3801\ : GlobalMux
    port map (
            O => \N__25800\,
            I => clk_12mhz
        );

    \I__3800\ : IoInMux
    port map (
            O => \N__25797\,
            I => \N__25794\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__25794\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25783\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25780\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25777\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25774\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25780\,
            I => \N__25771\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25777\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__3791\ : Odrv4
    port map (
            O => \N__25774\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__25771\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25759\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25756\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25753\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25759\,
            I => \N__25748\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__25756\,
            I => \N__25748\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25744\
        );

    \I__3783\ : Span4Mux_h
    port map (
            O => \N__25748\,
            I => \N__25741\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25738\
        );

    \I__3781\ : Span4Mux_h
    port map (
            O => \N__25744\,
            I => \N__25731\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__25741\,
            I => \N__25731\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25738\,
            I => \N__25731\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__25731\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25721\
        );

    \I__3775\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25718\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__25721\,
            I => \N__25715\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__25718\,
            I => \N__25709\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__25715\,
            I => \N__25709\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25706\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__25709\,
            I => \N__25703\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25706\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__25703\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25692\
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__25697\,
            I => \N__25689\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25686\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25683\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25692\,
            I => \N__25680\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25677\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25674\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25683\,
            I => \N__25671\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__25680\,
            I => \N__25666\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25666\
        );

    \I__3757\ : Span4Mux_h
    port map (
            O => \N__25674\,
            I => \N__25663\
        );

    \I__3756\ : Span12Mux_h
    port map (
            O => \N__25671\,
            I => \N__25660\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__25666\,
            I => \N__25657\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__25663\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__25660\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__25657\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25650\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25647\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25644\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25641\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__25638\,
            I => \N__25635\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25632\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25629\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25626\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25623\,
            I => \bfn_9_21_0_\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25620\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__3740\ : InMux
    port map (
            O => \N__25617\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__3737\ : Odrv12
    port map (
            O => \N__25608\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__3736\ : InMux
    port map (
            O => \N__25605\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25602\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25599\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25596\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25593\,
            I => \N__25590\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__25587\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25584\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25581\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__3727\ : InMux
    port map (
            O => \N__25578\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__3726\ : InMux
    port map (
            O => \N__25575\,
            I => \bfn_9_20_0_\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25572\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__25569\,
            I => \N__25566\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25562\
        );

    \I__3722\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25559\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25562\,
            I => \N__25556\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25553\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__25556\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__25553\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25541\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25538\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25535\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__25538\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__25535\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__3711\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__25527\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25524\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25521\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25515\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25512\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__25509\,
            I => \N__25506\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3701\ : Odrv12
    port map (
            O => \N__25500\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25497\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25494\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__3698\ : InMux
    port map (
            O => \N__25491\,
            I => \bfn_9_19_0_\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__25488\,
            I => \N__25485\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25482\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3693\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__25473\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__25464\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__3688\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__25458\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__3686\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__25449\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__25443\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3680\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__25428\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__25413\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__25401\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__25389\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__25383\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25374\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25374\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25374\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25365\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25365\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__25365\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25358\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25354\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25351\
        );

    \I__3652\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25347\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25342\
        );

    \I__3650\ : Span4Mux_v
    port map (
            O => \N__25351\,
            I => \N__25342\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25339\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25336\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__25342\,
            I => \N__25333\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25330\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__25336\,
            I => \N__25327\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__25333\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__3643\ : Odrv12
    port map (
            O => \N__25330\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__25327\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25317\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25313\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25309\
        );

    \I__3638\ : Span4Mux_v
    port map (
            O => \N__25313\,
            I => \N__25306\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25303\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25309\,
            I => \N__25296\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__25306\,
            I => \N__25296\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__25303\,
            I => \N__25296\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__25296\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__3632\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25287\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25287\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25287\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__25284\,
            I => \N__25280\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25275\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25275\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__25275\,
            I => \N__25272\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__25272\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__25266\,
            I => \N__25261\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25258\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25255\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__25261\,
            I => \N__25250\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25250\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25255\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__25250\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__3616\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25241\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25237\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__25241\,
            I => \N__25234\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25231\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25227\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__25234\,
            I => \N__25224\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__25231\,
            I => \N__25221\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25230\,
            I => \N__25218\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__25227\,
            I => \N__25213\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__25224\,
            I => \N__25213\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__25221\,
            I => \N__25208\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__25218\,
            I => \N__25208\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__25213\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__25208\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25200\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__25200\,
            I => \N__25196\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25192\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__25196\,
            I => \N__25189\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25186\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__25192\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__25189\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__25186\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25175\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25170\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__25175\,
            I => \N__25167\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25174\,
            I => \N__25164\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__25173\,
            I => \N__25161\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__25170\,
            I => \N__25156\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__25167\,
            I => \N__25156\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__25164\,
            I => \N__25153\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25150\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__25156\,
            I => \N__25147\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__25153\,
            I => \N__25144\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25141\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__25147\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__3581\ : Odrv4
    port map (
            O => \N__25144\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__25141\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__3579\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25131\,
            I => \N__25126\
        );

    \I__3577\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25123\
        );

    \I__3576\ : InMux
    port map (
            O => \N__25129\,
            I => \N__25120\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__25126\,
            I => \N__25114\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__25123\,
            I => \N__25114\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25120\,
            I => \N__25111\
        );

    \I__3572\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25108\
        );

    \I__3571\ : Span4Mux_v
    port map (
            O => \N__25114\,
            I => \N__25105\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__25111\,
            I => \N__25102\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__25108\,
            I => \N__25099\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__25105\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__25102\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__25099\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__3565\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25088\
        );

    \I__3564\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25084\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__25088\,
            I => \N__25081\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25078\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25084\,
            I => \N__25073\
        );

    \I__3560\ : Span4Mux_h
    port map (
            O => \N__25081\,
            I => \N__25073\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__25078\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__25073\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__3557\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__25060\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25057\
        );

    \I__3554\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25054\
        );

    \I__3553\ : Span12Mux_h
    port map (
            O => \N__25060\,
            I => \N__25051\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__25057\,
            I => \N__25048\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__25054\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__3550\ : Odrv12
    port map (
            O => \N__25051\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__25048\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__3548\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25037\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25034\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__25037\,
            I => \N__25029\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__25034\,
            I => \N__25026\
        );

    \I__3544\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25023\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25020\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__25029\,
            I => \N__25017\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__25026\,
            I => \N__25012\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25012\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25020\,
            I => \N__25009\
        );

    \I__3538\ : Span4Mux_v
    port map (
            O => \N__25017\,
            I => \N__25006\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__25012\,
            I => \N__25001\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__25009\,
            I => \N__25001\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__25006\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__25001\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24992\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24988\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24992\,
            I => \N__24985\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24982\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24979\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__24985\,
            I => \N__24974\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24982\,
            I => \N__24974\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24979\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__24974\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24960\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24957\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24954\
        );

    \I__3520\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24951\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__24960\,
            I => \N__24946\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24957\,
            I => \N__24946\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__24954\,
            I => \N__24943\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24951\,
            I => \N__24940\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__24946\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__24943\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__24940\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24929\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24925\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24929\,
            I => \N__24922\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24919\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24925\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3507\ : Odrv12
    port map (
            O => \N__24922\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24919\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24907\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24904\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24901\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24907\,
            I => \N__24893\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24893\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24901\,
            I => \N__24893\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24890\
        );

    \I__3498\ : Span4Mux_h
    port map (
            O => \N__24893\,
            I => \N__24885\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24885\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__24885\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24877\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24874\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24871\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24877\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24874\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24871\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24859\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24855\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24852\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24859\,
            I => \N__24849\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24846\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24855\,
            I => \N__24843\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24852\,
            I => \N__24840\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__24849\,
            I => \N__24835\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24846\,
            I => \N__24835\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__24843\,
            I => \N__24830\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__24840\,
            I => \N__24830\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__24835\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__24830\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24821\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24817\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__24821\,
            I => \N__24814\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24811\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24817\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__24814\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__24811\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24796\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24793\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24790\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__24796\,
            I => \N__24786\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__24793\,
            I => \N__24783\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24790\,
            I => \N__24780\
        );

    \I__3462\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24777\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__24786\,
            I => \N__24774\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__24783\,
            I => \N__24769\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__24780\,
            I => \N__24769\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24777\,
            I => \N__24766\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__24774\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__24769\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__3455\ : Odrv12
    port map (
            O => \N__24766\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24755\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24752\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24748\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24745\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24742\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__24748\,
            I => \N__24737\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__24745\,
            I => \N__24737\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24742\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24737\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24728\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24725\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24722\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24716\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__24722\,
            I => \N__24716\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24713\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__24716\,
            I => \N__24709\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24713\,
            I => \N__24706\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24703\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__24709\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__24706\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24703\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__24696\,
            I => \N__24693\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24689\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24686\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24689\,
            I => \N__24681\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__24686\,
            I => \N__24678\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24675\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24672\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__24681\,
            I => \N__24669\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__24678\,
            I => \N__24664\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24664\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24672\,
            I => \N__24661\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__24669\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24664\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__24661\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24649\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24646\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24643\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24649\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24646\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24643\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24631\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24628\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24625\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24622\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24617\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__24625\,
            I => \N__24617\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__24622\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__24617\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24607\
        );

    \I__3404\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24604\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24601\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__24607\,
            I => \N__24597\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__24604\,
            I => \N__24594\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24591\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24588\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__24597\,
            I => \N__24585\
        );

    \I__3397\ : Span12Mux_h
    port map (
            O => \N__24594\,
            I => \N__24578\
        );

    \I__3396\ : Span12Mux_s4_v
    port map (
            O => \N__24591\,
            I => \N__24578\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24578\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__24585\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__3393\ : Odrv12
    port map (
            O => \N__24578\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24573\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24570\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24567\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24564\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24561\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24558\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__24552\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24543\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__3381\ : InMux
    port map (
            O => \N__24540\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24537\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24531\,
            I => \N__24528\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__24528\,
            I => \N__24525\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__24525\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__3375\ : InMux
    port map (
            O => \N__24522\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__3373\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__24513\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24510\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__3370\ : InMux
    port map (
            O => \N__24507\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__24504\,
            I => \N__24501\
        );

    \I__3368\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24498\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24495\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24492\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24489\,
            I => \bfn_8_20_0_\
        );

    \I__3363\ : InMux
    port map (
            O => \N__24486\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24480\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24480\,
            I => \N__24477\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__24477\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24474\,
            I => \bfn_8_18_0_\
        );

    \I__3358\ : InMux
    port map (
            O => \N__24471\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__3357\ : InMux
    port map (
            O => \N__24468\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24465\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__3355\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__3353\ : Odrv12
    port map (
            O => \N__24456\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__3352\ : InMux
    port map (
            O => \N__24453\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24450\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__3350\ : InMux
    port map (
            O => \N__24447\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__24444\,
            I => \N__24441\
        );

    \I__3348\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24435\
        );

    \I__3346\ : Odrv12
    port map (
            O => \N__24435\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__3345\ : InMux
    port map (
            O => \N__24432\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24429\,
            I => \bfn_8_19_0_\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__24426\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24420\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__3340\ : InMux
    port map (
            O => \N__24417\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24414\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24411\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__24402\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24399\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24390\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24387\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__3329\ : InMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24381\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__3327\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__24375\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24364\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24361\
        );

    \I__3322\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24358\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24364\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__24361\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__24358\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24351\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24340\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24337\
        );

    \I__3314\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24334\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__24340\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__24337\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24334\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24327\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__3308\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24316\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24313\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24310\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24316\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24313\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__24310\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24303\,
            I => \bfn_8_12_0_\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24295\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24292\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24289\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__24295\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24292\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24289\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3295\ : InMux
    port map (
            O => \N__24282\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24271\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24268\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24265\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__24271\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24268\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24265\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3287\ : InMux
    port map (
            O => \N__24258\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__24255\,
            I => \N__24250\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__24254\,
            I => \N__24247\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24244\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24239\
        );

    \I__3282\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24239\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24244\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24239\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24234\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24227\
        );

    \I__3277\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24224\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__24227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24224\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24219\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24194\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24194\
        );

    \I__3271\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24194\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24194\
        );

    \I__3269\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24185\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24185\
        );

    \I__3267\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24185\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24185\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24180\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24180\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24155\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24155\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24155\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24155\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24152\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24149\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24180\,
            I => \N__24146\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24137\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24137\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24137\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24137\
        );

    \I__3252\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24128\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24128\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24128\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24128\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24119\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24119\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24119\
        );

    \I__3245\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24119\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24110\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24110\
        );

    \I__3242\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24110\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24110\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24155\,
            I => \N__24107\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__24152\,
            I => \N__24096\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__24149\,
            I => \N__24096\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__24146\,
            I => \N__24096\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24096\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24096\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24119\,
            I => \N__24091\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24091\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__24107\,
            I => \N__24088\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__24096\,
            I => \N__24085\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__24091\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__24088\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__24085\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24078\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__3226\ : InMux
    port map (
            O => \N__24075\,
            I => \N__24071\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24068\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__24071\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__24068\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3222\ : CEMux
    port map (
            O => \N__24063\,
            I => \N__24057\
        );

    \I__3221\ : CEMux
    port map (
            O => \N__24062\,
            I => \N__24054\
        );

    \I__3220\ : CEMux
    port map (
            O => \N__24061\,
            I => \N__24051\
        );

    \I__3219\ : CEMux
    port map (
            O => \N__24060\,
            I => \N__24048\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24045\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24042\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24039\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24036\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__24045\,
            I => \N__24033\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__24042\,
            I => \N__24026\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__24039\,
            I => \N__24026\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__24036\,
            I => \N__24026\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__24033\,
            I => \delay_measurement_inst.delay_tr_timer.N_344_i\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__24026\,
            I => \delay_measurement_inst.delay_tr_timer.N_344_i\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24013\
        );

    \I__3206\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24010\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24007\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__24013\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__24010\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__24007\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24000\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23989\
        );

    \I__3198\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23986\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23983\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23989\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23986\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__23983\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23976\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__23973\,
            I => \N__23970\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23965\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23962\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23959\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__23965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__23962\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23959\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23952\,
            I => \bfn_8_11_0_\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__23949\,
            I => \N__23946\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23941\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23938\
        );

    \I__3181\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23935\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23941\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23938\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23935\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23928\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__23925\,
            I => \N__23922\
        );

    \I__3175\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23917\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23914\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23911\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23917\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23914\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23911\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23904\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__23901\,
            I => \N__23898\
        );

    \I__3167\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23893\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23890\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23887\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23893\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23890\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23880\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23869\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23866\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23863\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23869\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__23866\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23856\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23845\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23842\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23839\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23845\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23842\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23839\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23832\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__23829\,
            I => \N__23826\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23821\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23818\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23815\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__23821\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23818\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23815\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23808\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__23805\,
            I => \N__23802\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23797\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23794\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23791\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23797\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23794\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23791\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23784\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23773\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23770\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23767\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23773\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__23770\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__23767\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23760\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23749\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23746\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23743\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23749\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__23746\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23743\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23736\,
            I => \bfn_8_10_0_\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23725\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23722\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23719\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23725\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23722\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23719\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23712\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23701\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23698\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23695\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23701\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23698\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23695\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23688\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23677\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23674\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23671\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23677\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23674\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23671\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23664\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23653\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23650\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23647\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__23653\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23650\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23647\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23640\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23629\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23626\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23623\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__23629\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23626\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23623\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23616\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23610\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23604\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23604\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23597\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__23600\,
            I => \N__23594\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23597\,
            I => \N__23590\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23587\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23584\
        );

    \I__3063\ : Odrv12
    port map (
            O => \N__23590\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23587\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__23584\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23577\,
            I => \bfn_8_9_0_\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23569\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23566\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23563\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23569\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23566\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__23563\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23556\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__23553\,
            I => \N__23550\
        );

    \I__3051\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23545\
        );

    \I__3050\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23542\
        );

    \I__3049\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23539\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__23545\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23542\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__23539\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23532\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__23529\,
            I => \N__23524\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__23528\,
            I => \N__23521\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23518\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23513\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23513\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23518\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__23513\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23508\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23497\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23494\
        );

    \I__3033\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23491\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__23497\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__23494\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23491\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23484\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__23481\,
            I => \N__23478\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23475\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23472\
        );

    \I__3025\ : Span4Mux_h
    port map (
            O => \N__23472\,
            I => \N__23469\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__23469\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__3023\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23463\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__23460\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23454\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23451\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__23451\,
            I => \N__23448\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__23448\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23442\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23439\
        );

    \I__3014\ : Span12Mux_v
    port map (
            O => \N__23439\,
            I => \N__23436\
        );

    \I__3013\ : Odrv12
    port map (
            O => \N__23436\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23427\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__23424\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__3006\ : Odrv12
    port map (
            O => \N__23415\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__23403\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__23400\,
            I => \N__23397\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__2998\ : Span12Mux_s7_h
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__2997\ : Odrv12
    port map (
            O => \N__23388\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__2993\ : Odrv12
    port map (
            O => \N__23376\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2992\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__23364\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23358\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__23355\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23349\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__23343\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2981\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23337\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__23334\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__23331\,
            I => \N__23328\
        );

    \I__2977\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__23325\,
            I => \N__23322\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__23319\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2973\ : InMux
    port map (
            O => \N__23316\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23313\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23310\,
            I => \bfn_7_13_0_\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23307\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23304\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23301\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23298\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__2966\ : CEMux
    port map (
            O => \N__23295\,
            I => \N__23290\
        );

    \I__2965\ : CEMux
    port map (
            O => \N__23294\,
            I => \N__23287\
        );

    \I__2964\ : CEMux
    port map (
            O => \N__23293\,
            I => \N__23284\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23290\,
            I => \N__23276\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23276\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__23284\,
            I => \N__23273\
        );

    \I__2960\ : CEMux
    port map (
            O => \N__23283\,
            I => \N__23270\
        );

    \I__2959\ : CEMux
    port map (
            O => \N__23282\,
            I => \N__23267\
        );

    \I__2958\ : CEMux
    port map (
            O => \N__23281\,
            I => \N__23264\
        );

    \I__2957\ : Span4Mux_v
    port map (
            O => \N__23276\,
            I => \N__23261\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__23273\,
            I => \N__23256\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23256\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23251\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__23264\,
            I => \N__23251\
        );

    \I__2952\ : Span4Mux_h
    port map (
            O => \N__23261\,
            I => \N__23246\
        );

    \I__2951\ : Span4Mux_h
    port map (
            O => \N__23256\,
            I => \N__23246\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__23251\,
            I => \N__23243\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__23246\,
            I => \delay_measurement_inst.delay_tr_timer.N_343_i\
        );

    \I__2948\ : Odrv4
    port map (
            O => \N__23243\,
            I => \delay_measurement_inst.delay_tr_timer.N_343_i\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__23232\,
            I => \N__23229\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__23229\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2943\ : InMux
    port map (
            O => \N__23226\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__2942\ : InMux
    port map (
            O => \N__23223\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23220\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23217\,
            I => \bfn_7_12_0_\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23214\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23211\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23208\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23205\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23202\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23199\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23196\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23193\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23190\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23187\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23184\,
            I => \bfn_7_11_0_\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23181\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23178\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23175\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23172\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__2924\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23166\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__23166\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__23163\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__23160\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__23157\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23151\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__23151\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__2917\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23145\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__23145\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23139\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23139\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__2913\ : InMux
    port map (
            O => \N__23136\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23133\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__23130\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23124\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__23124\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23118\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__23118\,
            I => \N__23115\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__23115\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__2905\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23109\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23106\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__23106\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23100\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__23100\,
            I => \N__23097\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__23097\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23091\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23087\
        );

    \I__2897\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23084\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__23087\,
            I => \N__23081\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23084\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__23081\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__23073\,
            I => \N__23069\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23066\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__23069\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__23066\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2888\ : InMux
    port map (
            O => \N__23061\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2887\ : InMux
    port map (
            O => \N__23058\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2886\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23050\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23047\
        );

    \I__2884\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23044\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23041\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23038\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23028\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__23041\,
            I => \N__23023\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23023\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23020\
        );

    \I__2877\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23011\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23011\
        );

    \I__2875\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23011\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23011\
        );

    \I__2873\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23006\
        );

    \I__2872\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23006\
        );

    \I__2871\ : Span4Mux_v
    port map (
            O => \N__23028\,
            I => \N__22999\
        );

    \I__2870\ : Span4Mux_v
    port map (
            O => \N__23023\,
            I => \N__22999\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__23020\,
            I => \N__22999\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__23011\,
            I => \N__22996\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__22993\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__22999\,
            I => \N__22990\
        );

    \I__2865\ : Span12Mux_s3_h
    port map (
            O => \N__22996\,
            I => \N__22985\
        );

    \I__2864\ : Sp12to4
    port map (
            O => \N__22993\,
            I => \N__22985\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__22990\,
            I => \N__22982\
        );

    \I__2862\ : Span12Mux_v
    port map (
            O => \N__22985\,
            I => \N__22979\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__22982\,
            I => \N__22976\
        );

    \I__2860\ : Odrv12
    port map (
            O => \N__22979\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__22976\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22968\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__22968\,
            I => \N__22965\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__22965\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__22959\,
            I => \N__22956\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__22956\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__22947\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22941\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__2847\ : Odrv12
    port map (
            O => \N__22938\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__22929\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22923\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22920\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__22920\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22914\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__22911\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22904\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22901\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22904\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__22901\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22896\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22889\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22886\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22889\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__22886\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22881\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22872\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__22872\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22865\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22865\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22862\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22857\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22848\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22848\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__22845\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22842\,
            I => \bfn_5_18_0_\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22833\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22833\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__22830\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22827\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__22818\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22808\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22805\
        );

    \I__2803\ : Span4Mux_h
    port map (
            O => \N__22808\,
            I => \N__22802\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22805\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__22802\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22797\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22787\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22784\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__22787\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22784\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22779\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22772\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__22775\,
            I => \N__22769\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22766\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22763\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__22766\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22763\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22758\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22752\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__22752\,
            I => \N__22748\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22745\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__22748\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22745\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22740\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22730\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__22733\,
            I => \N__22727\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22724\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22721\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__22724\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__22721\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22716\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22704\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22709\,
            I => \N__22704\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22704\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22701\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__22695\,
            I => \N__22692\
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__22692\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2764\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22683\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22683\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22683\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22680\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22674\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22670\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22667\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__22670\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22667\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22662\,
            I => \bfn_5_17_0_\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22649\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22646\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__22649\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22646\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22641\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22631\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22628\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__22631\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22628\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22623\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22616\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \N__22613\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22616\,
            I => \N__22610\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22607\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__22610\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__22607\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22602\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22593\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22593\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__22590\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22587\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__22578\,
            I => \N__22574\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22571\
        );

    \I__2725\ : Span4Mux_v
    port map (
            O => \N__22574\,
            I => \N__22565\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22565\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22562\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__22565\,
            I => \N__22559\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22556\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__2719\ : Span12Mux_s5_h
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__22553\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2717\ : Odrv12
    port map (
            O => \N__22550\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22545\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__22542\,
            I => \N__22538\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22535\
        );

    \I__2713\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22528\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22525\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22522\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__22528\,
            I => \N__22519\
        );

    \I__2708\ : Span4Mux_s3_h
    port map (
            O => \N__22525\,
            I => \N__22514\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22514\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__22519\,
            I => \N__22511\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__22514\,
            I => \N__22508\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__22511\,
            I => \N__22505\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__22508\,
            I => \N__22502\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__22505\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2700\ : InMux
    port map (
            O => \N__22497\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22491\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22486\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22483\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22480\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__22486\,
            I => \N__22475\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22475\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22472\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__22475\,
            I => \N__22469\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__22472\,
            I => \N__22466\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__22469\,
            I => \N__22463\
        );

    \I__2689\ : Sp12to4
    port map (
            O => \N__22466\,
            I => \N__22460\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__22463\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2687\ : Odrv12
    port map (
            O => \N__22460\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22455\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22444\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22441\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22438\
        );

    \I__2681\ : Sp12to4
    port map (
            O => \N__22444\,
            I => \N__22431\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22431\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22431\
        );

    \I__2678\ : Span12Mux_v
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__2677\ : Odrv12
    port map (
            O => \N__22428\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22425\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2675\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22417\
        );

    \I__2674\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22414\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \N__22411\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22408\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22402\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__22408\,
            I => \N__22397\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__22405\,
            I => \N__22397\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__22402\,
            I => \N__22394\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__22397\,
            I => \N__22391\
        );

    \I__2665\ : Span12Mux_s5_h
    port map (
            O => \N__22394\,
            I => \N__22388\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__22391\,
            I => \N__22385\
        );

    \I__2663\ : Odrv12
    port map (
            O => \N__22388\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__22385\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22380\,
            I => \bfn_5_16_0_\
        );

    \I__2660\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22373\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22370\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22373\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__22370\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22365\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22358\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22355\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22358\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__22355\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22350\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2650\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22340\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22337\
        );

    \I__2647\ : Odrv12
    port map (
            O => \N__22340\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22337\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22332\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2644\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22323\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22316\
        );

    \I__2642\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22316\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22316\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__22323\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__22316\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__22305\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22299\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22299\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__22296\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__22287\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__22284\,
            I => \N__22276\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \N__22273\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22270\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22267\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22256\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22256\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22256\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22256\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22256\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22267\,
            I => \N__22252\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__22256\,
            I => \N__22249\
        );

    \I__2618\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22246\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__22252\,
            I => \N__22243\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__22249\,
            I => \N__22238\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22238\
        );

    \I__2614\ : Span4Mux_v
    port map (
            O => \N__22243\,
            I => \N__22233\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__22238\,
            I => \N__22233\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__22230\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22224\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22221\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__22221\,
            I => \N__22218\
        );

    \I__2607\ : Sp12to4
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__22215\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22212\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22205\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22202\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22205\,
            I => \N__22196\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22196\
        );

    \I__2600\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22193\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__22196\,
            I => \N__22190\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22187\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__22190\,
            I => \N__22184\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22181\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22178\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__22181\,
            I => \N__22175\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__22178\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__22175\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22170\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22161\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22158\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22155\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22152\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22161\,
            I => \N__22147\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__22158\,
            I => \N__22147\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__22155\,
            I => \N__22144\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22141\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__22147\,
            I => \N__22138\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__22144\,
            I => \N__22135\
        );

    \I__2580\ : Span12Mux_s5_h
    port map (
            O => \N__22141\,
            I => \N__22132\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__22138\,
            I => \N__22129\
        );

    \I__2578\ : Span4Mux_v
    port map (
            O => \N__22135\,
            I => \N__22126\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__22132\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__22129\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__22126\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22119\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22109\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22105\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__22109\,
            I => \N__22102\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22099\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22105\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__22102\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__22099\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22085\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22081\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__22085\,
            I => \N__22078\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22075\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__22081\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__22078\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__22075\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22060\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22057\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22054\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__22060\,
            I => \N__22051\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__22057\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22054\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__22051\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2549\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22041\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22036\
        );

    \I__2547\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22033\
        );

    \I__2546\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22030\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__22036\,
            I => \N__22027\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22033\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__22030\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__22027\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__22020\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2540\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22009\
        );

    \I__2538\ : InMux
    port map (
            O => \N__22013\,
            I => \N__22006\
        );

    \I__2537\ : InMux
    port map (
            O => \N__22012\,
            I => \N__22003\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__22009\,
            I => \N__22000\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__22006\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__22003\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__22000\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21990\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21979\
        );

    \I__2528\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21976\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21973\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__21979\,
            I => \N__21970\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__21976\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21973\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__21970\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__21963\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__2521\ : InMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21957\,
            I => \N__21952\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21949\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21946\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__21952\,
            I => \N__21943\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21949\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21946\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__21943\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21918\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21918\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21918\
        );

    \I__2510\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21918\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21913\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21913\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21904\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21904\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21904\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21904\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21918\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__21913\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__21904\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__2498\ : Span4Mux_h
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__21882\,
            I => \N__21879\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__21879\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__21876\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21867\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__21864\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21858\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__21855\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21849\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21843\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__21834\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21824\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21820\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__21824\,
            I => \N__21817\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21814\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__21820\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__21817\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21814\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21800\
        );

    \I__2468\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21796\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__21800\,
            I => \N__21793\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21790\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21796\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__21793\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21790\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21775\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21772\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21769\
        );

    \I__2458\ : Span4Mux_v
    port map (
            O => \N__21775\,
            I => \N__21766\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21772\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21769\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__21766\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21756\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21756\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21753\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2451\ : IoInMux
    port map (
            O => \N__21750\,
            I => \N__21747\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21744\
        );

    \I__2449\ : Span12Mux_s1_v
    port map (
            O => \N__21744\,
            I => \N__21741\
        );

    \I__2448\ : Span12Mux_h
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__2447\ : Span12Mux_v
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2446\ : Odrv12
    port map (
            O => \N__21735\,
            I => pwm_output_c
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__21732\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__21729\,
            I => \N__21726\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21723\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__21720\,
            I => \N__21717\
        );

    \I__2440\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21714\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21714\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21705\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21705\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21694\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21677\
        );

    \I__2434\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21677\
        );

    \I__2433\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21677\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21677\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21677\
        );

    \I__2430\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21677\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21677\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21677\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__21694\,
            I => \N__21672\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21672\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__21669\,
            I => \N__21666\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__21666\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21657\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21657\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21646\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21629\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21629\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21629\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21629\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21629\
        );

    \I__2414\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21629\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21629\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21629\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__21646\,
            I => \N__21626\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21623\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__21626\,
            I => \N__21620\
        );

    \I__2408\ : Span12Mux_v
    port map (
            O => \N__21623\,
            I => \N__21617\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__21620\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__21617\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__21612\,
            I => \N__21608\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21583\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21583\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__21607\,
            I => \N__21579\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__21606\,
            I => \N__21575\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__21605\,
            I => \N__21571\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__21604\,
            I => \N__21567\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__21603\,
            I => \N__21559\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21541\
        );

    \I__2396\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21541\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21541\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21541\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21541\
        );

    \I__2392\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21541\
        );

    \I__2391\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21541\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21541\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21526\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21526\
        );

    \I__2387\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21526\
        );

    \I__2386\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21526\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21526\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21526\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21526\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21523\
        );

    \I__2381\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21506\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21506\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21506\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21506\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21506\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21506\
        );

    \I__2375\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21506\
        );

    \I__2374\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21506\
        );

    \I__2373\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21501\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21501\
        );

    \I__2371\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21494\
        );

    \I__2370\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21494\
        );

    \I__2369\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21494\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21491\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21488\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21485\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21482\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__21523\,
            I => \N__21477\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21477\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21472\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21472\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21463\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21463\
        );

    \I__2358\ : Sp12to4
    port map (
            O => \N__21485\,
            I => \N__21463\
        );

    \I__2357\ : Sp12to4
    port map (
            O => \N__21482\,
            I => \N__21463\
        );

    \I__2356\ : Span4Mux_h
    port map (
            O => \N__21477\,
            I => \N__21460\
        );

    \I__2355\ : Sp12to4
    port map (
            O => \N__21472\,
            I => \N__21455\
        );

    \I__2354\ : Span12Mux_v
    port map (
            O => \N__21463\,
            I => \N__21455\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__21460\,
            I => \N_19_1\
        );

    \I__2352\ : Odrv12
    port map (
            O => \N__21455\,
            I => \N_19_1\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21447\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__21447\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__2348\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__21438\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21432\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__21432\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__21429\,
            I => \N__21426\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__21423\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21417\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__21414\,
            I => \N__21411\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21408\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21405\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__21405\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21399\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__21390\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21384\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__21384\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__21381\,
            I => \N__21378\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21375\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__21369\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21360\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21360\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21354\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21348\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__21339\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21333\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21330\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21327\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21324\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21321\,
            I => \bfn_3_19_0_\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21318\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21312\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21312\,
            I => \N__21309\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__21309\,
            I => \N__21306\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__21306\,
            I => \N__21303\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__21303\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21294\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21291\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__21291\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21285\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21285\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__21282\,
            I => \N__21279\
        );

    \I__2294\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21276\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__21276\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21270\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__21270\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21261\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__21261\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__21255\,
            I => \N__21250\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21247\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21244\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__21250\,
            I => \N__21239\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21239\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__21244\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__21239\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__2278\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__21228\,
            I => \N__21224\
        );

    \I__2276\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21221\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__21224\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21221\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__2273\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__21213\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21203\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21199\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__21203\,
            I => \N__21196\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21193\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21199\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__21196\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__21193\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__2263\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__21180\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21171\,
            I => \N__21167\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21164\
        );

    \I__2256\ : Span4Mux_h
    port map (
            O => \N__21167\,
            I => \N__21161\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21158\
        );

    \I__2254\ : Sp12to4
    port map (
            O => \N__21161\,
            I => \N__21155\
        );

    \I__2253\ : Span4Mux_v
    port map (
            O => \N__21158\,
            I => \N__21152\
        );

    \I__2252\ : Odrv12
    port map (
            O => \N__21155\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__21152\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21144\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__21135\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21128\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21125\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21128\,
            I => \N__21122\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21119\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__21122\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__21119\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__21114\,
            I => \N__21107\
        );

    \I__2238\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21104\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__21112\,
            I => \N__21100\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__21111\,
            I => \N__21092\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21088\
        );

    \I__2234\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21085\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21082\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21077\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21077\
        );

    \I__2230\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21070\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21070\
        );

    \I__2228\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21070\
        );

    \I__2227\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21061\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21061\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21061\
        );

    \I__2224\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21061\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21054\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21054\
        );

    \I__2221\ : Span4Mux_s3_h
    port map (
            O => \N__21082\,
            I => \N__21054\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__21077\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__21070\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21061\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__21054\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__2216\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21041\
        );

    \I__2215\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21037\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__21041\,
            I => \N__21034\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21031\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21037\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__21034\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__21031\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__2209\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__21021\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__2207\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21011\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21001\
        );

    \I__2205\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21001\
        );

    \I__2204\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21001\
        );

    \I__2203\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21001\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__20998\
        );

    \I__2201\ : InMux
    port map (
            O => \N__21010\,
            I => \N__20995\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__21001\,
            I => \N__20988\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__20998\,
            I => \N__20988\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20995\,
            I => \N__20985\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20980\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20980\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__20988\,
            I => \N__20977\
        );

    \I__2194\ : Span4Mux_s3_h
    port map (
            O => \N__20985\,
            I => \N__20974\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__20980\,
            I => \N__20971\
        );

    \I__2192\ : Span12Mux_s3_h
    port map (
            O => \N__20977\,
            I => \N__20964\
        );

    \I__2191\ : Sp12to4
    port map (
            O => \N__20974\,
            I => \N__20964\
        );

    \I__2190\ : Sp12to4
    port map (
            O => \N__20971\,
            I => \N__20964\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__20964\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20961\,
            I => \bfn_3_18_0_\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20958\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20955\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20952\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20949\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__20940\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__20931\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20928\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20922\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20922\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20919\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20913\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20913\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20910\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__20901\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20892\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20889\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20883\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20883\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20880\,
            I => \bfn_3_16_0_\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20874\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__20868\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__20856\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20853\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20844\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20838\,
            I => \N__20833\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20828\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20828\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__20833\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20828\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20819\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20816\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20813\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20810\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__20813\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__20810\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20802\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__20793\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20784\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20784\,
            I => \N__20780\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20776\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__20780\,
            I => \N__20773\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20770\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20776\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__20773\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__20770\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20759\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20756\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20750\
        );

    \I__2118\ : Odrv12
    port map (
            O => \N__20753\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__20750\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20742\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__20742\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20739\,
            I => \N__20736\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20733\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__20724\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20718\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20718\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20715\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20706\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20706\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20703\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20697\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20694\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__20685\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20678\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20675\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20678\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20675\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20662\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20659\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20656\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20653\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20650\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__20656\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__20653\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__20650\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20638\
        );

    \I__2081\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20635\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20632\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20629\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__20635\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20632\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__20629\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20618\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20615\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20618\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20615\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20601\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__20601\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20595\,
            I => \N__20592\
        );

    \I__2065\ : Odrv12
    port map (
            O => \N__20592\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__2064\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20585\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20582\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20585\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__20582\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__20577\,
            I => \N__20574\
        );

    \I__2059\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20570\
        );

    \I__2058\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20566\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__20570\,
            I => \N__20563\
        );

    \I__2056\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20560\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__20566\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__20563\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20560\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2052\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20550\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__20550\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20543\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20539\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__20543\,
            I => \N__20536\
        );

    \I__2047\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20539\,
            I => pwm_duty_input_3
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__20536\,
            I => pwm_duty_input_3
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20533\,
            I => pwm_duty_input_3
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20520\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20512\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20509\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20506\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__20512\,
            I => \N__20503\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20498\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20498\
        );

    \I__2034\ : Span4Mux_s1_h
    port map (
            O => \N__20503\,
            I => \N__20495\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__20498\,
            I => pwm_duty_input_4
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20495\,
            I => pwm_duty_input_4
        );

    \I__2031\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20487\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20481\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20481\,
            I => \N__20478\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__20478\,
            I => \N__20475\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__20475\,
            I => \N__20472\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__20472\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__20469\,
            I => \N__20466\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20460\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__20454\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20448\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20448\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20445\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__2014\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__20433\,
            I => \N__20430\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__20427\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20421\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20421\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__2007\ : InMux
    port map (
            O => \N__20418\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__20415\,
            I => \N__20412\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20409\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20406\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__20400\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20394\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20394\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20391\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__20388\,
            I => \N__20385\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__20379\,
            I => \N__20376\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__20376\,
            I => \N__20373\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__20373\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__1991\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20367\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20364\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__20364\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20361\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20352\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__1983\ : Span4Mux_v
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__20343\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__20334\,
            I => \N__20331\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__20331\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20328\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20322\
        );

    \I__1975\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20316\
        );

    \I__1973\ : Span12Mux_v
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__1972\ : Odrv12
    port map (
            O => \N__20313\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__20304\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20301\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__1967\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20294\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20291\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__20294\,
            I => \N__20286\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20286\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__20286\,
            I => \N__20277\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20270\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20270\
        );

    \I__1960\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20270\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20263\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20263\
        );

    \I__1957\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20263\
        );

    \I__1956\ : Span4Mux_v
    port map (
            O => \N__20277\,
            I => \N__20256\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20256\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20256\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__20250\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__1949\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20241\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__20232\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20220\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__20220\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__20217\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20211\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__20208\,
            I => \N__20205\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__20205\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20199\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__20199\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__1933\ : InMux
    port map (
            O => \N__20196\,
            I => \bfn_2_17_0_\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__20181\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__20178\,
            I => \N__20175\
        );

    \I__1926\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__20169\,
            I => \N__20166\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__20166\,
            I => \N__20163\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__20163\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__20157\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20154\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__20145\,
            I => \N__20142\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__20139\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__20136\,
            I => \N__20133\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__20130\,
            I => \N__20127\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__1909\ : Span4Mux_s3_h
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__20118\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20112\
        );

    \I__1905\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20109\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__20109\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20106\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__1902\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20100\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__20100\,
            I => \N__20097\
        );

    \I__1900\ : Span12Mux_h
    port map (
            O => \N__20097\,
            I => \N__20094\
        );

    \I__1899\ : Odrv12
    port map (
            O => \N__20094\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__20091\,
            I => \N__20088\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20085\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__20085\,
            I => \N__20082\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__20082\,
            I => \N__20079\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__20076\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20070\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__20070\,
            I => \N__20067\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__20067\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__1889\ : InMux
    port map (
            O => \N__20064\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__1888\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20058\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__20058\,
            I => \N__20055\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__20049\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \N__20043\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__20031\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__20028\,
            I => \N__20025\
        );

    \I__1876\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__20019\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20016\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__1872\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__1869\ : Sp12to4
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__20001\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19989\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__19989\,
            I => \N__19986\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__19983\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__1861\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__19974\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__1858\ : InMux
    port map (
            O => \N__19971\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19965\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__1855\ : Span4Mux_s3_h
    port map (
            O => \N__19962\,
            I => \N__19959\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__19953\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__19935\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19926\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19923\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19920\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19914\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__19911\,
            I => \N__19908\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__19908\,
            I => \N__19905\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__19905\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__19902\,
            I => \N__19899\
        );

    \I__1834\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19896\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__19893\,
            I => \N__19890\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__19890\,
            I => \N__19887\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__19884\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19878\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19875\,
            I => \bfn_2_16_0_\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19872\,
            I => \bfn_2_14_0_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19869\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19866\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19863\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__19848\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__19833\,
            I => \N__19830\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__19827\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__19821\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__19806\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__19794\,
            I => \N__19791\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__19788\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__19779\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19776\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__1790\ : Span12Mux_h
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__1789\ : Odrv12
    port map (
            O => \N__19764\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__1787\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19755\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19746\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__19740\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__19734\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__1776\ : Span4Mux_v
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__19719\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19713\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19713\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__1771\ : InMux
    port map (
            O => \N__19710\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19703\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19700\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19697\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__19700\,
            I => \N__19694\
        );

    \I__1766\ : Span4Mux_h
    port map (
            O => \N__19697\,
            I => \N__19689\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__19694\,
            I => \N__19689\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__19686\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19683\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19680\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19677\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19674\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19671\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__19668\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19662\,
            I => \N__19659\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19659\,
            I => \N__19655\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__19655\,
            I => \current_shift_inst.PI_CTRL.N_306\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19652\,
            I => \current_shift_inst.PI_CTRL.N_306\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19641\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__19635\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19629\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__19629\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__19620\,
            I => \N__19617\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__19614\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19608\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__19608\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19602\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19602\,
            I => \N__19599\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__19596\,
            I => \N__19593\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__19593\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__19587\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19581\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19581\,
            I => \N__19578\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__19575\,
            I => \N__19572\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__19572\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__19566\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__1720\ : Span4Mux_h
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__19551\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1717\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__19545\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__19530\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__19524\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__1706\ : Span12Mux_v
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__19512\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19506\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19493\
        );

    \I__1700\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19493\
        );

    \I__1699\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19490\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19493\,
            I => pwm_duty_input_8
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__19490\,
            I => pwm_duty_input_8
        );

    \I__1696\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19478\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19478\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19475\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__19478\,
            I => \N__19472\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19469\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__19472\,
            I => pwm_duty_input_9
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__19469\,
            I => pwm_duty_input_9
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__19464\,
            I => \N__19460\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19456\
        );

    \I__1687\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19451\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19451\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19456\,
            I => \N__19448\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__19451\,
            I => pwm_duty_input_7
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__19448\,
            I => pwm_duty_input_7
        );

    \I__1682\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19436\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19436\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19433\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__19436\,
            I => pwm_duty_input_6
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__19433\,
            I => pwm_duty_input_6
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__19428\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__1676\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19417\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19412\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19412\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__19417\,
            I => \N__19409\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__19412\,
            I => pwm_duty_input_5
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__19409\,
            I => pwm_duty_input_5
        );

    \I__1669\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19400\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19397\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__19400\,
            I => \N__19392\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19397\,
            I => \N__19392\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__19392\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19380\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19380\
        );

    \I__1662\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19380\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__19380\,
            I => \current_shift_inst.PI_CTRL.N_120\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__19377\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19370\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19367\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__19370\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__19367\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19358\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19355\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__19358\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__19355\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19344\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1648\ : InMux
    port map (
            O => \N__19341\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19334\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19331\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19328\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__19331\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__19328\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__19317\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__1639\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__19311\,
            I => \N_6_0\
        );

    \I__1637\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__19305\,
            I => m38
        );

    \I__1635\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19298\
        );

    \I__1634\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19295\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19292\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__19295\,
            I => pwm_duty_input_0
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__19292\,
            I => pwm_duty_input_0
        );

    \I__1630\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19283\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19280\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__19283\,
            I => \N__19277\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__19280\,
            I => pwm_duty_input_1
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__19277\,
            I => pwm_duty_input_1
        );

    \I__1625\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19268\
        );

    \I__1624\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19265\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19262\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__19265\,
            I => pwm_duty_input_2
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__19262\,
            I => pwm_duty_input_2
        );

    \I__1620\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19254\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19251\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__1617\ : Span4Mux_v
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__19245\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1615\ : InMux
    port map (
            O => \N__19242\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__1614\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__19227\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19224\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__19209\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19206\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__1602\ : InMux
    port map (
            O => \N__19203\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__1601\ : InMux
    port map (
            O => \N__19200\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19197\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__1599\ : InMux
    port map (
            O => \N__19194\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__1598\ : InMux
    port map (
            O => \N__19191\,
            I => \bfn_1_17_0_\
        );

    \I__1597\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__19185\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__19182\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__1594\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__19176\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__1592\ : IoInMux
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__1590\ : IoSpan4Mux
    port map (
            O => \N__19167\,
            I => \N__19164\
        );

    \I__1589\ : IoSpan4Mux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__19161\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \I__1587\ : IoInMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19152\
        );

    \I__1585\ : Span4Mux_s3_v
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__19149\,
            I => \N__19146\
        );

    \I__1583\ : Sp12to4
    port map (
            O => \N__19146\,
            I => \N__19143\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__19137\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_14_21_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19158\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19173\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \phase_controller_inst2.stoper_tr.un1_start_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29912\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \current_shift_inst.timer_s1.running_RNI8ENL_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__38658\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_339_i_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__47166\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__49882\,
            CLKHFEN => \N__49884\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__49883\,
            RGB2PWM => \N__19314\,
            RGB1 => rgb_g_wire,
            CURREN => \N__49814\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19308\,
            RGB0PWM => \N__50418\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__23055\,
            in1 => \N__22281\,
            in2 => \N__22420\,
            in3 => \N__21018\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50915\,
            ce => 'H',
            sr => \N__50338\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21315\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50914\,
            ce => 'H',
            sr => \N__50345\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19388\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21897\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50914\,
            ce => 'H',
            sr => \N__50345\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22227\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50914\,
            ce => 'H',
            sr => \N__50345\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19179\,
            in2 => \_gnd_net_\,
            in3 => \N__19387\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50914\,
            ce => 'H',
            sr => \N__50345\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__21016\,
            in1 => \N__23036\,
            in2 => \N__22284\,
            in3 => \N__22452\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__22164\,
            in1 => \N__19188\,
            in2 => \N__19665\,
            in3 => \N__22280\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__21015\,
            in1 => \N__23035\,
            in2 => \N__22283\,
            in3 => \N__22494\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__23033\,
            in1 => \N__22279\,
            in2 => \N__22584\,
            in3 => \N__21017\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__21014\,
            in1 => \N__23034\,
            in2 => \N__22282\,
            in3 => \N__22541\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__22209\,
            in1 => \N__19404\,
            in2 => \_gnd_net_\,
            in3 => \N__19374\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50913\,
            ce => 'H',
            sr => \N__50352\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__22167\,
            in1 => \N__19362\,
            in2 => \N__23054\,
            in3 => \N__21010\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22165\,
            in2 => \_gnd_net_\,
            in3 => \N__22201\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__23037\,
            in1 => \N__19658\,
            in2 => \N__19182\,
            in3 => \N__22255\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23053\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50905\,
            ce => 'H',
            sr => \N__50374\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21206\,
            in2 => \_gnd_net_\,
            in3 => \N__21170\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21227\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20621\,
            in2 => \_gnd_net_\,
            in3 => \N__20642\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20665\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20681\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20588\,
            in2 => \_gnd_net_\,
            in3 => \N__20573\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19706\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19257\,
            in2 => \_gnd_net_\,
            in3 => \N__19242\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19239\,
            in2 => \_gnd_net_\,
            in3 => \N__19224\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19221\,
            in2 => \_gnd_net_\,
            in3 => \N__19206\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19824\,
            in2 => \_gnd_net_\,
            in3 => \N__19203\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49785\,
            in2 => \N__19785\,
            in3 => \N__19200\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20160\,
            in2 => \N__49815\,
            in3 => \N__19197\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49789\,
            in2 => \N__20115\,
            in3 => \N__19194\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20073\,
            in2 => \_gnd_net_\,
            in3 => \N__19191\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20028\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19980\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19881\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20451\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20424\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20397\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20370\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20340\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20310\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20229\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19341\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19338\,
            in1 => \N__20298\,
            in2 => \_gnd_net_\,
            in3 => \N__21558\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__19337\,
            in1 => \N__20297\,
            in2 => \N__21603\,
            in3 => \N__19323\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.m5_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__50417\,
            in1 => \N__43689\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.m38_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__50416\,
            in1 => \N__43688\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => m38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19301\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19459\,
            in2 => \_gnd_net_\,
            in3 => \N__19420\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19499\,
            in1 => \N__19484\,
            in2 => \N__19503\,
            in3 => \N__19442\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19500\,
            in1 => \N__19485\,
            in2 => \N__19464\,
            in3 => \N__19443\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20546\,
            in1 => \N__20516\,
            in2 => \N__19428\,
            in3 => \N__19421\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19373\,
            in1 => \N__19403\,
            in2 => \N__19350\,
            in3 => \N__22208\,
            lcout => \current_shift_inst.PI_CTRL.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__22489\,
            in1 => \N__22447\,
            in2 => \N__22542\,
            in3 => \N__20490\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__20993\,
            in1 => \N__23032\,
            in2 => \N__19377\,
            in3 => \N__22166\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__23031\,
            in1 => \N__20994\,
            in2 => \_gnd_net_\,
            in3 => \N__19361\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22531\,
            in2 => \_gnd_net_\,
            in3 => \N__22422\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22448\,
            in1 => \N__22490\,
            in2 => \N__19668\,
            in3 => \N__22577\,
            lcout => \current_shift_inst.PI_CTRL.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__19647\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19611\,
            in2 => \_gnd_net_\,
            in3 => \N__19626\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19590\,
            in2 => \_gnd_net_\,
            in3 => \N__19605\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19569\,
            in2 => \_gnd_net_\,
            in3 => \N__19584\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19548\,
            in2 => \_gnd_net_\,
            in3 => \N__19563\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19527\,
            in2 => \_gnd_net_\,
            in3 => \N__19542\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19509\,
            in2 => \_gnd_net_\,
            in3 => \N__19521\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19773\,
            in1 => \_gnd_net_\,
            in2 => \N__19761\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19737\,
            in2 => \_gnd_net_\,
            in3 => \N__19752\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19716\,
            in2 => \_gnd_net_\,
            in3 => \N__19731\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \_gnd_net_\,
            in3 => \N__19710\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21113\,
            in1 => \N__19707\,
            in2 => \_gnd_net_\,
            in3 => \N__19683\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21040\,
            in2 => \_gnd_net_\,
            in3 => \N__19680\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21254\,
            in2 => \_gnd_net_\,
            in3 => \N__19677\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20666\,
            in2 => \_gnd_net_\,
            in3 => \N__19674\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20779\,
            in2 => \_gnd_net_\,
            in3 => \N__19671\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20836\,
            in2 => \_gnd_net_\,
            in3 => \N__19872\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20569\,
            in2 => \_gnd_net_\,
            in3 => \N__19869\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20641\,
            in2 => \_gnd_net_\,
            in3 => \N__19866\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19863\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20837\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21044\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20762\,
            in2 => \_gnd_net_\,
            in3 => \N__20783\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19860\,
            in2 => \N__19845\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19818\,
            in2 => \N__19803\,
            in3 => \N__19776\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20193\,
            in2 => \N__20178\,
            in3 => \N__20154\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20151\,
            in2 => \N__20136\,
            in3 => \N__20106\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20103\,
            in2 => \N__20091\,
            in3 => \N__20064\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20061\,
            in2 => \N__20046\,
            in3 => \N__20016\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20013\,
            in2 => \N__19998\,
            in3 => \N__19971\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19968\,
            in2 => \N__19950\,
            in3 => \N__19920\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19917\,
            in2 => \N__19902\,
            in3 => \N__19875\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20484\,
            in2 => \N__20469\,
            in3 => \N__20445\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20280\,
            in2 => \N__20442\,
            in3 => \N__20418\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20283\,
            in2 => \N__20415\,
            in3 => \N__20391\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20281\,
            in2 => \N__20388\,
            in3 => \N__20361\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20284\,
            in2 => \N__20358\,
            in3 => \N__20328\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20282\,
            in2 => \N__20325\,
            in3 => \N__20301\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20285\,
            in2 => \N__20247\,
            in3 => \N__20217\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20214\,
            in1 => \N__20202\,
            in2 => \_gnd_net_\,
            in3 => \N__20196\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20691\,
            in1 => \N__20682\,
            in2 => \N__20670\,
            in3 => \N__21097\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20643\,
            in1 => \N__20622\,
            in2 => \N__20610\,
            in3 => \N__21099\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20598\,
            in1 => \N__20589\,
            in2 => \N__20577\,
            in3 => \N__21098\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__20553\,
            in1 => \N__20547\,
            in2 => \N__20526\,
            in3 => \N__20515\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22421\,
            in2 => \_gnd_net_\,
            in3 => \N__22570\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21700\,
            in1 => \N__21652\,
            in2 => \N__21605\,
            in3 => \N__20700\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21651\,
            in1 => \N__21574\,
            in2 => \N__20712\,
            in3 => \N__21699\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__21698\,
            in1 => \N__20721\,
            in2 => \N__21604\,
            in3 => \N__21650\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__21656\,
            in1 => \N__21582\,
            in2 => \N__20898\,
            in3 => \N__21704\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__21703\,
            in1 => \N__21655\,
            in2 => \N__21607\,
            in3 => \N__20916\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21653\,
            in1 => \N__21578\,
            in2 => \N__20937\,
            in3 => \N__21701\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21702\,
            in1 => \N__21654\,
            in2 => \N__21606\,
            in3 => \N__20925\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21649\,
            in1 => \N__21570\,
            in2 => \N__20739\,
            in3 => \N__21697\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21147\,
            in2 => \N__21114\,
            in3 => \N__21110\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20730\,
            in2 => \_gnd_net_\,
            in3 => \N__20715\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21024\,
            in2 => \_gnd_net_\,
            in3 => \N__20703\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21216\,
            in2 => \_gnd_net_\,
            in3 => \N__20694\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20946\,
            in2 => \_gnd_net_\,
            in3 => \N__20928\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20745\,
            in2 => \_gnd_net_\,
            in3 => \N__20919\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20805\,
            in2 => \_gnd_net_\,
            in3 => \N__20910\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20907\,
            in2 => \_gnd_net_\,
            in3 => \N__20889\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20886\,
            in2 => \_gnd_net_\,
            in3 => \N__20880\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__20877\,
            in1 => \N__21103\,
            in2 => \N__20865\,
            in3 => \N__20853\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__20850\,
            in1 => \N__20841\,
            in2 => \N__21112\,
            in3 => \N__20823\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__20799\,
            in2 => \N__20790\,
            in3 => \N__20763\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21267\,
            in1 => \N__21258\,
            in2 => \N__21234\,
            in3 => \N__21095\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21210\,
            in1 => \N__21186\,
            in2 => \N__21177\,
            in3 => \N__21091\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__21141\,
            in1 => \N__21132\,
            in2 => \N__21111\,
            in3 => \N__21045\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21435\,
            in1 => \N__21852\,
            in2 => \N__21873\,
            in3 => \N__21861\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21933\,
            in1 => \N__22088\,
            in2 => \_gnd_net_\,
            in3 => \N__20961\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_1_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21927\,
            in1 => \N__22013\,
            in2 => \_gnd_net_\,
            in3 => \N__20958\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_2_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21934\,
            in1 => \N__22112\,
            in2 => \_gnd_net_\,
            in3 => \N__20955\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_3_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__22040\,
            in2 => \_gnd_net_\,
            in3 => \N__20952\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_4_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21935\,
            in1 => \N__22064\,
            in2 => \_gnd_net_\,
            in3 => \N__20949\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_5_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21929\,
            in1 => \N__21955\,
            in2 => \_gnd_net_\,
            in3 => \N__21330\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_6_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21936\,
            in1 => \N__21983\,
            in2 => \_gnd_net_\,
            in3 => \N__21327\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_7_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21930\,
            in1 => \N__21779\,
            in2 => \_gnd_net_\,
            in3 => \N__21324\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__50821\,
            ce => 'H',
            sr => \N__50389\
        );

    \pwm_generator_inst.counter_8_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__21803\,
            in2 => \_gnd_net_\,
            in3 => \N__21321\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__50811\,
            ce => 'H',
            sr => \N__50393\
        );

    \pwm_generator_inst.counter_9_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21827\,
            in1 => \N__21931\,
            in2 => \_gnd_net_\,
            in3 => \N__21318\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50811\,
            ce => 'H',
            sr => \N__50393\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__22329\,
            in1 => \N__31311\,
            in2 => \_gnd_net_\,
            in3 => \N__28628\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50894\,
            ce => 'H',
            sr => \N__50358\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30696\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50877\,
            ce => 'H',
            sr => \N__50369\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21288\,
            in2 => \N__21300\,
            in3 => \N__22092\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21273\,
            in2 => \N__21282\,
            in3 => \N__22017\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21420\,
            in2 => \N__21429\,
            in3 => \N__22116\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21402\,
            in2 => \N__21414\,
            in3 => \N__22044\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21387\,
            in2 => \N__21396\,
            in3 => \N__22068\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21372\,
            in2 => \N__21381\,
            in3 => \N__21960\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21357\,
            in2 => \N__21366\,
            in3 => \N__21987\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21351\,
            in2 => \N__21345\,
            in3 => \N__21783\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21336\,
            in2 => \N__21720\,
            in3 => \N__21807\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21759\,
            in2 => \N__21444\,
            in3 => \N__21831\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21753\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50854\,
            ce => 'H',
            sr => \N__50375\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22815\,
            in1 => \N__22677\,
            in2 => \N__22659\,
            in3 => \N__23076\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22343\,
            in2 => \_gnd_net_\,
            in3 => \N__22377\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22362\,
            in1 => \N__22794\,
            in2 => \N__21732\,
            in3 => \N__21840\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__21662\,
            in1 => \N__21611\,
            in2 => \N__21729\,
            in3 => \N__21710\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21711\,
            in1 => \N__21663\,
            in2 => \N__21612\,
            in3 => \N__21450\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22751\,
            in1 => \N__22869\,
            in2 => \N__22733\,
            in3 => \N__22893\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22688\,
            in2 => \_gnd_net_\,
            in3 => \N__22709\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22854\,
            in1 => \N__22838\,
            in2 => \N__21876\,
            in3 => \N__22908\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22853\,
            in1 => \N__22839\,
            in2 => \N__22619\,
            in3 => \N__22634\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22689\,
            in1 => \N__22776\,
            in2 => \N__22713\,
            in3 => \N__22376\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22347\,
            in1 => \N__22361\,
            in2 => \N__21864\,
            in3 => \N__21846\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22907\,
            in2 => \_gnd_net_\,
            in3 => \N__22599\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22811\,
            in1 => \N__22790\,
            in2 => \N__21855\,
            in3 => \N__23072\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22652\,
            in2 => \_gnd_net_\,
            in3 => \N__22673\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22598\,
            in1 => \N__22868\,
            in2 => \N__22775\,
            in3 => \N__22892\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21823\,
            in1 => \N__21799\,
            in2 => \_gnd_net_\,
            in3 => \N__21778\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22108\,
            in2 => \_gnd_net_\,
            in3 => \N__22084\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__22063\,
            in1 => \N__22039\,
            in2 => \N__22020\,
            in3 => \N__22012\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__21982\,
            in2 => \N__21963\,
            in3 => \N__21956\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36869\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50803\,
            ce => 'H',
            sr => \N__50390\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23090\,
            in2 => \_gnd_net_\,
            in3 => \N__41795\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50795\,
            ce => 'H',
            sr => \N__50394\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25064\,
            in1 => \N__25041\,
            in2 => \_gnd_net_\,
            in3 => \N__32561\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50900\,
            ce => \N__31703\,
            sr => \N__50339\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23601\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50895\,
            ce => \N__23281\,
            sr => \N__50346\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22326\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__22328\,
            in1 => \_gnd_net_\,
            in2 => \N__28629\,
            in3 => \N__31310\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_344_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22327\,
            in2 => \_gnd_net_\,
            in3 => \N__28624\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_343_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37275\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50878\,
            ce => 'H',
            sr => \N__50359\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36578\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50855\,
            ce => 'H',
            sr => \N__50370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22755\,
            in1 => \N__22620\,
            in2 => \N__22737\,
            in3 => \N__22638\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22311\,
            in1 => \N__22302\,
            in2 => \N__22296\,
            in3 => \N__22293\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23094\,
            in2 => \N__41805\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23352\,
            in2 => \N__41703\,
            in3 => \N__22212\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23412\,
            in2 => \N__41631\,
            in3 => \N__22170\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50940\,
            in2 => \N__42669\,
            in3 => \N__22119\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42568\,
            in2 => \N__23400\,
            in3 => \N__22545\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23373\,
            in2 => \N__46899\,
            in3 => \N__22497\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46950\,
            in2 => \N__23481\,
            in3 => \N__22455\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38202\,
            in2 => \N__42462\,
            in3 => \N__22425\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__50835\,
            ce => 'H',
            sr => \N__50376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22962\,
            in2 => \N__42384\,
            in3 => \N__22380\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22971\,
            in2 => \N__42318\,
            in3 => \N__22365\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23457\,
            in2 => \N__42243\,
            in3 => \N__22350\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23421\,
            in2 => \N__46838\,
            in3 => \N__22332\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23445\,
            in2 => \N__46248\,
            in3 => \N__22740\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42984\,
            in2 => \N__23331\,
            in3 => \N__22716\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22944\,
            in2 => \N__42915\,
            in3 => \N__22701\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22698\,
            in2 => \N__42846\,
            in3 => \N__22680\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__50822\,
            ce => 'H',
            sr => \N__50380\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23361\,
            in2 => \N__42786\,
            in3 => \N__22662\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22926\,
            in2 => \N__42732\,
            in3 => \N__22641\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22935\,
            in2 => \N__43527\,
            in3 => \N__22623\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23238\,
            in2 => \N__43473\,
            in3 => \N__22602\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43413\,
            in2 => \N__23385\,
            in3 => \N__22587\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22953\,
            in2 => \N__43362\,
            in3 => \N__22896\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23112\,
            in2 => \N__43296\,
            in3 => \N__22881\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22878\,
            in2 => \N__43242\,
            in3 => \N__22857\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__50812\,
            ce => 'H',
            sr => \N__50383\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22917\,
            in2 => \N__43173\,
            in3 => \N__22842\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23433\,
            in2 => \N__43116\,
            in3 => \N__22827\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22824\,
            in2 => \N__43992\,
            in3 => \N__22797\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23121\,
            in2 => \N__43932\,
            in3 => \N__22779\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23103\,
            in2 => \N__43872\,
            in3 => \N__22758\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23340\,
            in2 => \N__43812\,
            in3 => \N__23061\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46608\,
            in1 => \N__23466\,
            in2 => \_gnd_net_\,
            in3 => \N__23058\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50804\,
            ce => 'H',
            sr => \N__50385\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36233\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36275\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36942\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36605\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37052\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36495\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50796\,
            ce => 'H',
            sr => \N__50388\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36821\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__50391\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37226\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__50391\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36899\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__50391\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37184\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__50391\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36014\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__50391\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25714\,
            in1 => \N__25698\,
            in2 => \_gnd_net_\,
            in3 => \N__32485\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32487\,
            in1 => \N__24610\,
            in2 => \_gnd_net_\,
            in3 => \N__24635\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25264\,
            in1 => \N__25240\,
            in2 => \_gnd_net_\,
            in3 => \N__32486\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32494\,
            in1 => \N__25906\,
            in2 => \_gnd_net_\,
            in3 => \N__25867\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50901\,
            ce => \N__32169\,
            sr => \N__50306\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28801\,
            in1 => \N__32493\,
            in2 => \_gnd_net_\,
            in3 => \N__28774\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26215\,
            in1 => \N__26245\,
            in2 => \_gnd_net_\,
            in3 => \N__32384\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32385\,
            in1 => \N__24932\,
            in2 => \_gnd_net_\,
            in3 => \N__24910\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26020\,
            in1 => \N__26050\,
            in2 => \_gnd_net_\,
            in3 => \N__32382\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32383\,
            in1 => \N__25316\,
            in2 => \_gnd_net_\,
            in3 => \N__25350\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25119\,
            in1 => \N__26158\,
            in2 => \N__25697\,
            in3 => \N__26095\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23607\,
            in1 => \N__23613\,
            in2 => \N__23130\,
            in3 => \N__23127\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26214\,
            in1 => \N__24789\,
            in2 => \N__32747\,
            in3 => \N__31801\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25230\,
            in2 => \_gnd_net_\,
            in3 => \N__28764\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25033\,
            in1 => \N__25063\,
            in2 => \_gnd_net_\,
            in3 => \N__32364\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31401\,
            in1 => \N__23142\,
            in2 => \_gnd_net_\,
            in3 => \N__26367\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__23169\,
            in2 => \N__23163\,
            in3 => \N__23148\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__24751\,
            in1 => \_gnd_net_\,
            in2 => \N__23160\,
            in3 => \N__24721\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24900\,
            in1 => \N__24862\,
            in2 => \N__25173\,
            in3 => \N__24963\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24684\,
            in1 => \N__25896\,
            in2 => \N__23157\,
            in3 => \N__23154\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24712\,
            in1 => \N__26011\,
            in2 => \N__25956\,
            in3 => \N__25747\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23574\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50879\,
            ce => \N__23282\,
            sr => \N__50332\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23548\,
            in2 => \N__23600\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23573\,
            in2 => \N__23528\,
            in3 => \N__23136\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23500\,
            in2 => \N__23553\,
            in3 => \N__23133\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23824\,
            in2 => \N__23529\,
            in3 => \N__23199\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23800\,
            in2 => \N__23505\,
            in3 => \N__23196\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23776\,
            in2 => \N__23829\,
            in3 => \N__23193\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23752\,
            in2 => \N__23805\,
            in3 => \N__23190\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23728\,
            in2 => \N__23781\,
            in3 => \N__23187\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50868\,
            ce => \N__23283\,
            sr => \N__50340\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23704\,
            in2 => \N__23757\,
            in3 => \N__23184\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23680\,
            in2 => \N__23733\,
            in3 => \N__23181\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23656\,
            in2 => \N__23709\,
            in3 => \N__23178\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23632\,
            in2 => \N__23685\,
            in3 => \N__23175\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24016\,
            in2 => \N__23661\,
            in3 => \N__23172\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23992\,
            in2 => \N__23637\,
            in3 => \N__23226\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23968\,
            in2 => \N__24021\,
            in3 => \N__23223\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23944\,
            in2 => \N__23997\,
            in3 => \N__23220\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50856\,
            ce => \N__23294\,
            sr => \N__50347\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23920\,
            in2 => \N__23973\,
            in3 => \N__23217\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23896\,
            in2 => \N__23949\,
            in3 => \N__23214\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23872\,
            in2 => \N__23925\,
            in3 => \N__23211\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23848\,
            in2 => \N__23901\,
            in3 => \N__23208\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24367\,
            in2 => \N__23877\,
            in3 => \N__23205\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24343\,
            in2 => \N__23853\,
            in3 => \N__23202\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24319\,
            in2 => \N__24372\,
            in3 => \N__23316\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24298\,
            in2 => \N__24348\,
            in3 => \N__23313\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50845\,
            ce => \N__23293\,
            sr => \N__50353\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24274\,
            in2 => \N__24324\,
            in3 => \N__23310\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50836\,
            ce => \N__23295\,
            sr => \N__50360\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24300\,
            in2 => \N__24254\,
            in3 => \N__23307\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50836\,
            ce => \N__23295\,
            sr => \N__50360\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24230\,
            in2 => \N__24279\,
            in3 => \N__23304\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50836\,
            ce => \N__23295\,
            sr => \N__50360\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24074\,
            in2 => \N__24255\,
            in3 => \N__23301\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50836\,
            ce => \N__23295\,
            sr => \N__50360\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23298\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50836\,
            ce => \N__23295\,
            sr => \N__50360\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36165\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50813\,
            ce => \N__36198\,
            sr => \N__50371\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37023\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50805\,
            ce => 'H',
            sr => \N__50373\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36725\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50805\,
            ce => 'H',
            sr => \N__50373\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36443\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50805\,
            ce => 'H',
            sr => \N__50373\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36399\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50797\,
            ce => 'H',
            sr => \N__50377\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36983\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50797\,
            ce => 'H',
            sr => \N__50377\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36362\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50797\,
            ce => 'H',
            sr => \N__50377\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36524\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50797\,
            ce => 'H',
            sr => \N__50377\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35966\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50787\,
            ce => 'H',
            sr => \N__50381\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37149\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50787\,
            ce => 'H',
            sr => \N__50381\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36648\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50787\,
            ce => 'H',
            sr => \N__50381\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36320\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50787\,
            ce => 'H',
            sr => \N__50381\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37101\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50787\,
            ce => 'H',
            sr => \N__50381\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33952\,
            in1 => \N__34339\,
            in2 => \N__35802\,
            in3 => \N__30329\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34338\,
            in1 => \N__33953\,
            in2 => \N__35886\,
            in3 => \N__33284\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36761\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50774\,
            ce => 'H',
            sr => \N__50386\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__41568\,
            in1 => \N__46329\,
            in2 => \_gnd_net_\,
            in3 => \N__46770\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50774\,
            ce => 'H',
            sr => \N__50386\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__46769\,
            in1 => \N__46607\,
            in2 => \N__46386\,
            in3 => \N__42519\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50774\,
            ce => 'H',
            sr => \N__50386\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36684\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50774\,
            ce => 'H',
            sr => \N__50386\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37316\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50774\,
            ce => 'H',
            sr => \N__50386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25786\,
            in1 => \N__25763\,
            in2 => \_gnd_net_\,
            in3 => \N__32492\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25199\,
            in1 => \N__25174\,
            in2 => \_gnd_net_\,
            in3 => \N__32489\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24824\,
            in1 => \N__24799\,
            in2 => \_gnd_net_\,
            in3 => \N__32491\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25871\,
            in1 => \N__25907\,
            in2 => \_gnd_net_\,
            in3 => \N__32490\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32488\,
            in1 => \N__28873\,
            in2 => \_gnd_net_\,
            in3 => \N__28847\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24612\,
            in1 => \N__24636\,
            in2 => \_gnd_net_\,
            in3 => \N__32433\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50887\,
            ce => \N__32074\,
            sr => \N__50307\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24928\,
            in1 => \N__24911\,
            in2 => \_gnd_net_\,
            in3 => \N__32432\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50887\,
            ce => \N__32074\,
            sr => \N__50307\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24654\,
            in1 => \N__24685\,
            in2 => \_gnd_net_\,
            in3 => \N__32390\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27341\,
            in1 => \N__27312\,
            in2 => \_gnd_net_\,
            in3 => \N__32388\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32389\,
            in1 => \N__24882\,
            in2 => \_gnd_net_\,
            in3 => \N__24858\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32812\,
            in1 => \N__32223\,
            in2 => \N__31745\,
            in3 => \N__25357\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32387\,
            in1 => \_gnd_net_\,
            in2 => \N__24995\,
            in3 => \N__24964\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25087\,
            in1 => \N__25129\,
            in2 => \_gnd_net_\,
            in3 => \N__32386\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25032\,
            in1 => \N__26609\,
            in2 => \N__27317\,
            in3 => \N__28839\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24213\,
            in1 => \N__23593\,
            in2 => \_gnd_net_\,
            in3 => \N__23577\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24209\,
            in1 => \N__23572\,
            in2 => \_gnd_net_\,
            in3 => \N__23556\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24214\,
            in1 => \N__23549\,
            in2 => \_gnd_net_\,
            in3 => \N__23532\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24210\,
            in1 => \N__23527\,
            in2 => \_gnd_net_\,
            in3 => \N__23508\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24215\,
            in1 => \N__23501\,
            in2 => \_gnd_net_\,
            in3 => \N__23484\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__23825\,
            in2 => \_gnd_net_\,
            in3 => \N__23808\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24216\,
            in1 => \N__23801\,
            in2 => \_gnd_net_\,
            in3 => \N__23784\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24212\,
            in1 => \N__23777\,
            in2 => \_gnd_net_\,
            in3 => \N__23760\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__50869\,
            ce => \N__24062\,
            sr => \N__50323\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24167\,
            in1 => \N__23753\,
            in2 => \_gnd_net_\,
            in3 => \N__23736\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24171\,
            in1 => \N__23729\,
            in2 => \_gnd_net_\,
            in3 => \N__23712\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24164\,
            in1 => \N__23705\,
            in2 => \_gnd_net_\,
            in3 => \N__23688\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24168\,
            in1 => \N__23681\,
            in2 => \_gnd_net_\,
            in3 => \N__23664\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24165\,
            in1 => \N__23657\,
            in2 => \_gnd_net_\,
            in3 => \N__23640\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24169\,
            in1 => \N__23633\,
            in2 => \_gnd_net_\,
            in3 => \N__23616\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24166\,
            in1 => \N__24017\,
            in2 => \_gnd_net_\,
            in3 => \N__24000\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24170\,
            in1 => \N__23993\,
            in2 => \_gnd_net_\,
            in3 => \N__23976\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__50857\,
            ce => \N__24060\,
            sr => \N__50333\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24172\,
            in1 => \N__23969\,
            in2 => \_gnd_net_\,
            in3 => \N__23952\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24176\,
            in1 => \N__23945\,
            in2 => \_gnd_net_\,
            in3 => \N__23928\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__23921\,
            in2 => \_gnd_net_\,
            in3 => \N__23904\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24177\,
            in1 => \N__23897\,
            in2 => \_gnd_net_\,
            in3 => \N__23880\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24174\,
            in1 => \N__23873\,
            in2 => \_gnd_net_\,
            in3 => \N__23856\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24178\,
            in1 => \N__23849\,
            in2 => \_gnd_net_\,
            in3 => \N__23832\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24175\,
            in1 => \N__24368\,
            in2 => \_gnd_net_\,
            in3 => \N__24351\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24179\,
            in1 => \N__24344\,
            in2 => \_gnd_net_\,
            in3 => \N__24327\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__50846\,
            ce => \N__24061\,
            sr => \N__50341\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24203\,
            in1 => \N__24320\,
            in2 => \_gnd_net_\,
            in3 => \N__24303\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24207\,
            in1 => \N__24299\,
            in2 => \_gnd_net_\,
            in3 => \N__24282\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24204\,
            in1 => \N__24275\,
            in2 => \_gnd_net_\,
            in3 => \N__24258\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24208\,
            in1 => \N__24253\,
            in2 => \_gnd_net_\,
            in3 => \N__24234\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24205\,
            in1 => \N__24231\,
            in2 => \_gnd_net_\,
            in3 => \N__24219\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24075\,
            in1 => \N__24206\,
            in2 => \_gnd_net_\,
            in3 => \N__24078\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50837\,
            ce => \N__24063\,
            sr => \N__50348\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31482\,
            lcout => \phase_controller_inst2.start_latched\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50823\,
            ce => 'H',
            sr => \N__50354\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34315\,
            in1 => \N__35534\,
            in2 => \N__33963\,
            in3 => \N__30407\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__38347\,
            in1 => \N__33859\,
            in2 => \N__38394\,
            in3 => \N__34316\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34198\,
            in1 => \N__33784\,
            in2 => \N__35937\,
            in3 => \N__33138\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33783\,
            in1 => \N__34197\,
            in2 => \N__35142\,
            in3 => \N__30065\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33781\,
            in1 => \N__34132\,
            in2 => \N__35196\,
            in3 => \N__30102\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34131\,
            in1 => \N__33018\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__49784\,
            in1 => \N__24384\,
            in2 => \_gnd_net_\,
            in3 => \N__31839\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34133\,
            in1 => \N__33782\,
            in2 => \N__38616\,
            in3 => \N__38571\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31869\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34130\,
            in2 => \N__24426\,
            in3 => \N__33017\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24423\,
            in2 => \N__25569\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29808\,
            in2 => \N__25398\,
            in3 => \N__28673\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28674\,
            in1 => \N__33484\,
            in2 => \N__25488\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25386\,
            in2 => \N__33670\,
            in3 => \N__24417\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33488\,
            in2 => \N__26514\,
            in3 => \N__24414\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33502\,
            in2 => \N__25410\,
            in3 => \N__24411\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33489\,
            in2 => \N__24408\,
            in3 => \N__24399\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33503\,
            in2 => \N__24396\,
            in3 => \N__24387\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24483\,
            in2 => \N__33762\,
            in3 => \N__24474\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33581\,
            in2 => \N__25440\,
            in3 => \N__24471\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25446\,
            in2 => \N__33763\,
            in3 => \N__24468\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33585\,
            in2 => \N__25479\,
            in3 => \N__24465\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24462\,
            in2 => \N__33764\,
            in3 => \N__24453\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33589\,
            in2 => \N__26481\,
            in3 => \N__24450\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25461\,
            in2 => \N__33765\,
            in3 => \N__24447\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33593\,
            in2 => \N__24444\,
            in3 => \N__24432\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33690\,
            in2 => \N__25425\,
            in3 => \N__24429\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25455\,
            in2 => \N__33867\,
            in3 => \N__24540\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33694\,
            in2 => \N__26451\,
            in3 => \N__24537\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24534\,
            in2 => \N__33868\,
            in3 => \N__24522\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33698\,
            in2 => \N__24519\,
            in3 => \N__24510\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26697\,
            in2 => \N__33869\,
            in3 => \N__24507\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33702\,
            in2 => \N__24504\,
            in3 => \N__24495\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25470\,
            in2 => \N__33870\,
            in3 => \N__24492\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33746\,
            in2 => \N__33321\,
            in3 => \N__24489\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26727\,
            in2 => \N__33896\,
            in3 => \N__24486\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33750\,
            in2 => \N__26886\,
            in3 => \N__24573\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26622\,
            in2 => \N__33897\,
            in3 => \N__24570\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33754\,
            in2 => \N__26652\,
            in3 => \N__24567\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24555\,
            in2 => \N__33898\,
            in3 => \N__24564\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33758\,
            in2 => \N__24549\,
            in3 => \N__24561\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__25815\,
            in2 => \N__34750\,
            in3 => \N__24558\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__36078\,
            in2 => \N__33971\,
            in3 => \N__30788\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__34333\,
            in1 => \N__30330\,
            in2 => \N__33970\,
            in3 => \N__35801\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__30612\,
            in1 => \N__33895\,
            in2 => \N__28694\,
            in3 => \N__34335\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24759\,
            in1 => \N__24732\,
            in2 => \_gnd_net_\,
            in3 => \N__32666\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50896\,
            ce => \N__31696\,
            sr => \N__50283\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32664\,
            in1 => \N__25265\,
            in2 => \_gnd_net_\,
            in3 => \N__25245\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50896\,
            ce => \N__31696\,
            sr => \N__50283\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24634\,
            in1 => \N__24611\,
            in2 => \_gnd_net_\,
            in3 => \N__32665\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50896\,
            ce => \N__31696\,
            sr => \N__50283\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32660\,
            in1 => \N__26109\,
            in2 => \_gnd_net_\,
            in3 => \N__26124\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50888\,
            ce => \N__31700\,
            sr => \N__50293\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24820\,
            in1 => \N__24804\,
            in2 => \_gnd_net_\,
            in3 => \N__32662\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50888\,
            ce => \N__31700\,
            sr => \N__50293\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25092\,
            in1 => \N__25134\,
            in2 => \_gnd_net_\,
            in3 => \N__32663\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50888\,
            ce => \N__31700\,
            sr => \N__50293\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25195\,
            in1 => \N__25179\,
            in2 => \_gnd_net_\,
            in3 => \N__32661\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50888\,
            ce => \N__31700\,
            sr => \N__50293\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25312\,
            in1 => \N__25362\,
            in2 => \_gnd_net_\,
            in3 => \N__32606\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26394\,
            in1 => \N__26373\,
            in2 => \_gnd_net_\,
            in3 => \N__32607\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32604\,
            in1 => \N__24692\,
            in2 => \_gnd_net_\,
            in3 => \N__24653\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24881\,
            in1 => \N__24864\,
            in2 => \_gnd_net_\,
            in3 => \N__32605\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32603\,
            in1 => \N__24933\,
            in2 => \_gnd_net_\,
            in3 => \N__24912\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24996\,
            in1 => \N__24969\,
            in2 => \_gnd_net_\,
            in3 => \N__32608\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50880\,
            ce => \N__31702\,
            sr => \N__50300\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24880\,
            in1 => \N__24863\,
            in2 => \_gnd_net_\,
            in3 => \N__32564\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50870\,
            ce => \N__32176\,
            sr => \N__50308\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32639\,
            in1 => \N__24825\,
            in2 => \_gnd_net_\,
            in3 => \N__24800\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50870\,
            ce => \N__32176\,
            sr => \N__50308\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31762\,
            in1 => \N__31740\,
            in2 => \_gnd_net_\,
            in3 => \N__32565\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50870\,
            ce => \N__32176\,
            sr => \N__50308\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32667\,
            in1 => \N__24758\,
            in2 => \_gnd_net_\,
            in3 => \N__24731\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27340\,
            in1 => \N__27316\,
            in2 => \_gnd_net_\,
            in3 => \N__32650\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32644\,
            in1 => \_gnd_net_\,
            in2 => \N__24696\,
            in3 => \N__24652\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28806\,
            in1 => \N__32648\,
            in2 => \_gnd_net_\,
            in3 => \N__28778\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25269\,
            in1 => \_gnd_net_\,
            in2 => \N__32694\,
            in3 => \N__25244\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25791\,
            in1 => \N__25762\,
            in2 => \_gnd_net_\,
            in3 => \N__32649\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50858\,
            ce => \N__32134\,
            sr => \N__50316\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25203\,
            in1 => \N__25178\,
            in2 => \_gnd_net_\,
            in3 => \N__32654\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32659\,
            in1 => \N__25130\,
            in2 => \_gnd_net_\,
            in3 => \N__25091\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32653\,
            in1 => \N__25068\,
            in2 => \_gnd_net_\,
            in3 => \N__25040\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24991\,
            in1 => \N__24965\,
            in2 => \_gnd_net_\,
            in3 => \N__32656\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32651\,
            in1 => \N__26250\,
            in2 => \_gnd_net_\,
            in3 => \N__26222\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28878\,
            in1 => \N__28846\,
            in2 => \_gnd_net_\,
            in3 => \N__32655\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32652\,
            in1 => \_gnd_net_\,
            in2 => \N__25728\,
            in3 => \N__25696\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50847\,
            ce => \N__32177\,
            sr => \N__50324\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__25380\,
            in1 => \N__28218\,
            in2 => \N__28247\,
            in3 => \N__25371\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32611\,
            in1 => \N__25991\,
            in2 => \_gnd_net_\,
            in3 => \N__25966\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__25379\,
            in1 => \N__28217\,
            in2 => \N__28248\,
            in3 => \N__25370\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26393\,
            in1 => \N__26368\,
            in2 => \_gnd_net_\,
            in3 => \N__32612\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__28322\,
            in1 => \N__25283\,
            in2 => \N__28350\,
            in3 => \N__25293\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25361\,
            in1 => \N__25320\,
            in2 => \_gnd_net_\,
            in3 => \N__32658\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50824\,
            ce => \N__32178\,
            sr => \N__50342\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__25292\,
            in1 => \N__28349\,
            in2 => \N__25284\,
            in3 => \N__28323\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32657\,
            in1 => \N__25987\,
            in2 => \_gnd_net_\,
            in3 => \N__25970\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50824\,
            ce => \N__32178\,
            sr => \N__50342\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26610\,
            in1 => \N__26319\,
            in2 => \_gnd_net_\,
            in3 => \N__32693\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50814\,
            ce => \N__31704\,
            sr => \N__50349\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34288\,
            in1 => \N__35094\,
            in2 => \N__33976\,
            in3 => \N__31910\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34289\,
            in1 => \N__35438\,
            in2 => \N__33977\,
            in3 => \N__30182\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33787\,
            in1 => \N__34247\,
            in2 => \N__35195\,
            in3 => \N__30101\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__49726\,
            in1 => \N__28672\,
            in2 => \_gnd_net_\,
            in3 => \N__25544\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__33785\,
            in1 => \N__34248\,
            in2 => \N__31917\,
            in3 => \N__35093\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34246\,
            in1 => \N__33786\,
            in2 => \N__35237\,
            in3 => \N__30134\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__29816\,
            in1 => \N__29772\,
            in2 => \N__29712\,
            in3 => \N__34245\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34177\,
            in1 => \N__35315\,
            in2 => \N__33855\,
            in3 => \N__32981\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36164\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50788\,
            ce => \N__36196\,
            sr => \N__50364\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__35351\,
            in1 => \N__34176\,
            in2 => \N__29688\,
            in3 => \N__33661\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34183\,
            in1 => \N__38064\,
            in2 => \N__33789\,
            in3 => \N__38031\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30372\,
            in1 => \N__33628\,
            in2 => \N__35748\,
            in3 => \N__34191\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__33627\,
            in1 => \N__38112\,
            in2 => \N__34287\,
            in3 => \N__30218\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__37940\,
            in1 => \N__33629\,
            in2 => \N__37983\,
            in3 => \N__34190\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34180\,
            in1 => \N__35316\,
            in2 => \N__33788\,
            in3 => \N__32988\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30027\,
            in1 => \N__33621\,
            in2 => \N__35058\,
            in3 => \N__34182\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__33626\,
            in1 => \N__30249\,
            in2 => \N__34286\,
            in3 => \N__35487\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__35238\,
            in1 => \N__33622\,
            in2 => \N__30138\,
            in3 => \N__34181\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25565\,
            in2 => \N__25548\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29809\,
            in2 => \N__29790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33490\,
            in2 => \N__26736\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25530\,
            in2 => \N__33671\,
            in3 => \N__25524\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33494\,
            in2 => \N__26706\,
            in3 => \N__25521\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25518\,
            in2 => \N__33672\,
            in3 => \N__25512\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33498\,
            in2 => \N__25509\,
            in3 => \N__25497\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26673\,
            in2 => \N__33673\,
            in3 => \N__25494\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33674\,
            in2 => \N__26634\,
            in3 => \N__25491\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25614\,
            in2 => \N__33863\,
            in3 => \N__25605\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33678\,
            in2 => \N__26466\,
            in3 => \N__25602\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26745\,
            in2 => \N__33864\,
            in3 => \N__25599\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33682\,
            in2 => \N__26811\,
            in3 => \N__25596\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25593\,
            in2 => \N__33865\,
            in3 => \N__25584\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33686\,
            in2 => \N__26895\,
            in3 => \N__25581\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26436\,
            in2 => \N__33866\,
            in3 => \N__25578\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33706\,
            in2 => \N__26496\,
            in3 => \N__25575\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26790\,
            in2 => \N__33871\,
            in3 => \N__25572\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33710\,
            in2 => \N__26904\,
            in3 => \N__25650\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26685\,
            in2 => \N__33872\,
            in3 => \N__25647\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33714\,
            in2 => \N__26802\,
            in3 => \N__25644\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26769\,
            in2 => \N__33873\,
            in3 => \N__25641\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33718\,
            in2 => \N__25638\,
            in3 => \N__25629\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26715\,
            in2 => \N__33874\,
            in3 => \N__25626\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33875\,
            in2 => \N__26919\,
            in3 => \N__25623\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26817\,
            in2 => \N__33967\,
            in3 => \N__25620\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33879\,
            in2 => \N__27006\,
            in3 => \N__25617\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26664\,
            in2 => \N__33968\,
            in3 => \N__25830\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33883\,
            in2 => \N__26874\,
            in3 => \N__25827\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27012\,
            in2 => \N__33969\,
            in3 => \N__25824\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33887\,
            in2 => \N__28644\,
            in3 => \N__25821\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33888\,
            in1 => \N__34336\,
            in2 => \_gnd_net_\,
            in3 => \N__25818\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25809\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_er_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29084\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50889\,
            ce => \N__26277\,
            sr => \N__50262\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25787\,
            in1 => \N__25764\,
            in2 => \_gnd_net_\,
            in3 => \N__32682\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50881\,
            ce => \N__31694\,
            sr => \N__50269\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32681\,
            in1 => \N__25724\,
            in2 => \_gnd_net_\,
            in3 => \N__25695\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50881\,
            ce => \N__31694\,
            sr => \N__50269\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25995\,
            in1 => \N__25971\,
            in2 => \_gnd_net_\,
            in3 => \N__32683\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50881\,
            ce => \N__31694\,
            sr => \N__50269\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__29300\,
            in1 => \N__25929\,
            in2 => \N__25920\,
            in3 => \N__29642\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__25928\,
            in1 => \N__29301\,
            in2 => \N__29643\,
            in3 => \N__25916\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26172\,
            in1 => \N__32679\,
            in2 => \_gnd_net_\,
            in3 => \N__26187\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50872\,
            ce => \N__31695\,
            sr => \N__50275\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32678\,
            in1 => \N__26057\,
            in2 => \_gnd_net_\,
            in3 => \N__26031\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50872\,
            ce => \N__31695\,
            sr => \N__50275\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25908\,
            in1 => \N__25872\,
            in2 => \_gnd_net_\,
            in3 => \N__32680\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50872\,
            ce => \N__31695\,
            sr => \N__50275\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__29351\,
            in1 => \N__25851\,
            in2 => \N__25842\,
            in3 => \N__29327\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__25850\,
            in1 => \N__29352\,
            in2 => \N__29328\,
            in3 => \N__25838\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32745\,
            in1 => \N__32768\,
            in2 => \_gnd_net_\,
            in3 => \N__32610\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50860\,
            ce => \N__31697\,
            sr => \N__50284\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32609\,
            in1 => \N__26246\,
            in2 => \_gnd_net_\,
            in3 => \N__26223\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50860\,
            ce => \N__31697\,
            sr => \N__50284\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__28272\,
            in1 => \N__28295\,
            in2 => \N__26136\,
            in3 => \N__26070\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26069\,
            in1 => \N__28271\,
            in2 => \N__28299\,
            in3 => \N__26132\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32674\,
            in1 => \N__26167\,
            in2 => \_gnd_net_\,
            in3 => \N__26183\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26168\,
            in1 => \_gnd_net_\,
            in2 => \N__26139\,
            in3 => \N__32676\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50849\,
            ce => \N__32171\,
            sr => \N__50294\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32673\,
            in1 => \N__26107\,
            in2 => \_gnd_net_\,
            in3 => \N__26120\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26108\,
            in1 => \_gnd_net_\,
            in2 => \N__26073\,
            in3 => \N__32675\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50849\,
            ce => \N__32171\,
            sr => \N__50294\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26061\,
            in1 => \N__26027\,
            in2 => \_gnd_net_\,
            in3 => \N__32677\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50849\,
            ce => \N__32171\,
            sr => \N__50294\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__28035\,
            in1 => \N__26304\,
            in2 => \N__28065\,
            in3 => \N__26295\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31810\,
            in1 => \N__31778\,
            in2 => \_gnd_net_\,
            in3 => \N__32670\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32672\,
            in1 => \_gnd_net_\,
            in2 => \N__26307\,
            in3 => \N__31811\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50838\,
            ce => \N__32133\,
            sr => \N__50301\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__28034\,
            in1 => \N__26303\,
            in2 => \N__28064\,
            in3 => \N__26294\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31741\,
            in1 => \N__31766\,
            in2 => \_gnd_net_\,
            in3 => \N__32671\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31224\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.start_latched\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50826\,
            ce => 'H',
            sr => \N__50309\
        );

    \phase_controller_inst1.stoper_tr.running_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__29074\,
            in1 => \N__26266\,
            in2 => \_gnd_net_\,
            in3 => \N__26286\,
            lcout => \phase_controller_inst1.running\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50826\,
            ce => 'H',
            sr => \N__50309\
        );

    \phase_controller_inst1.stoper_hc.m42_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101011101"
        )
    port map (
            in0 => \N__31223\,
            in1 => \N__29073\,
            in2 => \N__26268\,
            in3 => \N__27726\,
            lcout => \phase_controller_inst1.N_43\,
            ltout => \phase_controller_inst1.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_sbtinv_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26280\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.m41_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__31222\,
            in1 => \N__29072\,
            in2 => \N__26267\,
            in3 => \N__27725\,
            lcout => \phase_controller_inst1.N_42\,
            ltout => \phase_controller_inst1.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32172\,
            in2 => \N__26424\,
            in3 => \N__27707\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50826\,
            ce => 'H',
            sr => \N__50309\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010110010"
        )
    port map (
            in0 => \N__26418\,
            in1 => \N__28446\,
            in2 => \N__26409\,
            in3 => \N__28470\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31402\,
            in1 => \N__32622\,
            in2 => \_gnd_net_\,
            in3 => \N__31358\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32623\,
            in1 => \_gnd_net_\,
            in2 => \N__26421\,
            in3 => \N__31403\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50816\,
            ce => \N__32135\,
            sr => \N__50317\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__26417\,
            in1 => \N__28445\,
            in2 => \N__26408\,
            in3 => \N__28469\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__26562\,
            in1 => \N__28391\,
            in2 => \N__26546\,
            in3 => \N__28422\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__26571\,
            in1 => \N__28493\,
            in2 => \N__26331\,
            in3 => \N__28194\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100001101"
        )
    port map (
            in0 => \N__28193\,
            in1 => \N__26570\,
            in2 => \N__28497\,
            in3 => \N__26327\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26389\,
            in1 => \N__26369\,
            in2 => \_gnd_net_\,
            in3 => \N__32626\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50807\,
            ce => \N__32170\,
            sr => \N__50325\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32624\,
            in1 => \N__26604\,
            in2 => \_gnd_net_\,
            in3 => \N__26318\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26605\,
            in1 => \_gnd_net_\,
            in2 => \N__26574\,
            in3 => \N__32625\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50807\,
            ce => \N__32170\,
            sr => \N__50325\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__26561\,
            in1 => \N__28392\,
            in2 => \N__26547\,
            in3 => \N__28418\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34282\,
            in1 => \N__35273\,
            in2 => \N__33989\,
            in3 => \N__32924\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38517\,
            in1 => \N__35050\,
            in2 => \_gnd_net_\,
            in3 => \N__30016\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30183\,
            in1 => \N__33915\,
            in2 => \N__35439\,
            in3 => \N__34285\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34284\,
            in1 => \N__35483\,
            in2 => \N__33978\,
            in3 => \N__30247\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__35051\,
            in1 => \N__34283\,
            in2 => \N__30023\,
            in3 => \N__33911\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__33959\,
            in1 => \N__34213\,
            in2 => \N__30536\,
            in3 => \N__35393\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34212\,
            in1 => \N__33962\,
            in2 => \N__38355\,
            in3 => \N__38387\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38499\,
            in1 => \N__35344\,
            in2 => \_gnd_net_\,
            in3 => \N__29680\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__33960\,
            in1 => \N__33083\,
            in2 => \N__35844\,
            in3 => \N__34215\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38500\,
            in1 => \N__35224\,
            in2 => \_gnd_net_\,
            in3 => \N__30133\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33961\,
            in1 => \N__34214\,
            in2 => \N__35936\,
            in3 => \N__33137\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__38612\,
            in2 => \N__33981\,
            in3 => \N__38570\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__35574\,
            in1 => \N__34195\,
            in2 => \N__30288\,
            in3 => \N__33920\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34196\,
            in1 => \N__36125\,
            in2 => \N__33980\,
            in3 => \N__31109\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30064\,
            in1 => \N__33927\,
            in2 => \N__35138\,
            in3 => \N__34193\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34194\,
            in1 => \N__35573\,
            in2 => \N__33979\,
            in3 => \N__30283\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34179\,
            in1 => \N__38060\,
            in2 => \N__33916\,
            in3 => \N__38030\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33793\,
            in1 => \N__34178\,
            in2 => \N__35355\,
            in3 => \N__29684\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__38101\,
            in1 => \N__38528\,
            in2 => \_gnd_net_\,
            in3 => \N__30217\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38529\,
            in1 => \N__35791\,
            in2 => \_gnd_net_\,
            in3 => \N__30322\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38527\,
            in1 => \N__35482\,
            in2 => \_gnd_net_\,
            in3 => \N__30248\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38526\,
            in1 => \N__35182\,
            in2 => \_gnd_net_\,
            in3 => \N__30100\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30581\,
            in1 => \N__33935\,
            in2 => \N__35654\,
            in3 => \N__34244\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34243\,
            in1 => \N__35744\,
            in2 => \N__33983\,
            in3 => \N__30371\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38530\,
            in1 => \N__35131\,
            in2 => \_gnd_net_\,
            in3 => \N__30066\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34241\,
            in1 => \N__35274\,
            in2 => \N__33982\,
            in3 => \N__32931\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__30287\,
            in1 => \N__34240\,
            in2 => \_gnd_net_\,
            in3 => \N__35567\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35690\,
            in1 => \N__38532\,
            in2 => \_gnd_net_\,
            in3 => \N__33350\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__30414\,
            in1 => \N__33931\,
            in2 => \N__35538\,
            in3 => \N__34242\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35431\,
            in1 => \N__38531\,
            in2 => \_gnd_net_\,
            in3 => \N__30181\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__33285\,
            in1 => \N__33941\,
            in2 => \N__35882\,
            in3 => \N__34320\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34318\,
            in1 => \N__37982\,
            in2 => \N__33985\,
            in3 => \N__37944\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__26784\,
            in1 => \N__26775\,
            in2 => \_gnd_net_\,
            in3 => \N__34716\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__33937\,
            in1 => \N__35843\,
            in2 => \N__34341\,
            in3 => \N__33087\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__26763\,
            in1 => \N__26754\,
            in2 => \_gnd_net_\,
            in3 => \N__34717\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__34324\,
            in1 => \N__35694\,
            in2 => \N__33357\,
            in3 => \N__33945\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__35394\,
            in1 => \N__34319\,
            in2 => \N__30540\,
            in3 => \N__33936\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34317\,
            in1 => \N__38111\,
            in2 => \N__33984\,
            in3 => \N__30219\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33948\,
            in1 => \N__34326\,
            in2 => \N__35613\,
            in3 => \N__30896\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34327\,
            in1 => \N__33946\,
            in2 => \N__36126\,
            in3 => \N__31113\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__34704\,
            in1 => \N__26865\,
            in2 => \_gnd_net_\,
            in3 => \N__26859\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__26850\,
            in1 => \N__26838\,
            in2 => \_gnd_net_\,
            in3 => \N__34702\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34705\,
            in1 => \N__26832\,
            in2 => \_gnd_net_\,
            in3 => \N__26823\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__34325\,
            in1 => \N__33947\,
            in2 => \N__35658\,
            in3 => \N__30582\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__34703\,
            in1 => \_gnd_net_\,
            in2 => \N__27033\,
            in3 => \N__27021\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__33987\,
            in1 => \N__34329\,
            in2 => \N__30792\,
            in3 => \N__36077\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__34328\,
            in1 => \N__33988\,
            in2 => \N__30903\,
            in3 => \N__35612\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26997\,
            in2 => \N__26991\,
            in3 => \N__29008\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28977\,
            in1 => \N__26982\,
            in2 => \N__26976\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28941\,
            in1 => \N__26967\,
            in2 => \N__26958\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26949\,
            in2 => \N__26943\,
            in3 => \N__28923\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28905\,
            in1 => \N__26934\,
            in2 => \N__26928\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27180\,
            in2 => \N__27168\,
            in3 => \N__29277\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27159\,
            in2 => \N__28740\,
            in3 => \N__29256\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27153\,
            in2 => \N__27144\,
            in3 => \N__29235\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27135\,
            in2 => \N__27123\,
            in3 => \N__29214\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29196\,
            in1 => \N__27111\,
            in2 => \N__27099\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29178\,
            in1 => \N__27090\,
            in2 => \N__27078\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27069\,
            in2 => \N__27060\,
            in3 => \N__29160\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27051\,
            in2 => \N__27042\,
            in3 => \N__29142\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27252\,
            in2 => \N__27246\,
            in3 => \N__29445\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27234\,
            in2 => \N__27228\,
            in3 => \N__29427\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31638\,
            in2 => \N__31566\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28731\,
            in2 => \N__28725\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27219\,
            in2 => \N__27210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27201\,
            in2 => \N__27189\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29091\,
            in2 => \N__28887\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29019\,
            in2 => \N__28716\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27408\,
            in2 => \N__27387\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27375\,
            in2 => \N__27351\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.un4_running_cry_30_THRU_LUT4_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27411\,
            lcout => \phase_controller_inst2.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__29511\,
            in1 => \N__27398\,
            in2 => \N__29490\,
            in3 => \N__31347\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__31346\,
            in1 => \N__29489\,
            in2 => \N__27402\,
            in3 => \N__29510\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__27278\,
            in1 => \N__29846\,
            in2 => \N__27369\,
            in3 => \N__29465\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__29466\,
            in1 => \N__27365\,
            in2 => \N__29847\,
            in3 => \N__27279\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27342\,
            in1 => \N__27321\,
            in2 => \_gnd_net_\,
            in3 => \N__32640\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50839\,
            ce => \N__31698\,
            sr => \N__50285\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27270\,
            in2 => \N__27261\,
            in3 => \N__27703\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27561\,
            in2 => \N__27549\,
            in3 => \N__28011\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27540\,
            in2 => \N__27531\,
            in3 => \N__27978\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27522\,
            in2 => \N__27516\,
            in3 => \N__27960\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27507\,
            in2 => \N__27495\,
            in3 => \N__27942\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27924\,
            in1 => \N__27486\,
            in2 => \N__27477\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27465\,
            in2 => \N__27456\,
            in3 => \N__27906\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27447\,
            in2 => \N__27438\,
            in3 => \N__27888\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27429\,
            in2 => \N__27420\,
            in3 => \N__27870\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27687\,
            in2 => \N__27675\,
            in3 => \N__28173\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27666\,
            in2 => \N__27654\,
            in3 => \N__28155\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28137\,
            in1 => \N__27645\,
            in2 => \N__27636\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28119\,
            in1 => \N__27627\,
            in2 => \N__27615\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28101\,
            in1 => \N__32706\,
            in2 => \N__27603\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28083\,
            in1 => \N__27582\,
            in2 => \N__27594\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27576\,
            in2 => \N__27570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31491\,
            in2 => \N__31551\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27852\,
            in2 => \N__27840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27825\,
            in2 => \N__27813\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27798\,
            in2 => \N__27789\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27777\,
            in2 => \N__27771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27762\,
            in2 => \N__27756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27744\,
            in2 => \N__27738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un4_running_cry_30_THRU_LUT4_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27729\,
            lcout => \phase_controller_inst1.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27717\,
            in1 => \N__27708\,
            in2 => \N__27992\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.N_42_i\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32104\,
            in1 => \N__28010\,
            in2 => \_gnd_net_\,
            in3 => \N__27996\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32108\,
            in1 => \N__27977\,
            in2 => \N__27993\,
            in3 => \N__27963\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32105\,
            in1 => \N__27959\,
            in2 => \_gnd_net_\,
            in3 => \N__27945\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32109\,
            in1 => \N__27941\,
            in2 => \_gnd_net_\,
            in3 => \N__27927\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32106\,
            in1 => \N__27923\,
            in2 => \_gnd_net_\,
            in3 => \N__27909\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32110\,
            in1 => \N__27905\,
            in2 => \_gnd_net_\,
            in3 => \N__27891\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32107\,
            in1 => \N__27887\,
            in2 => \_gnd_net_\,
            in3 => \N__27873\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__50799\,
            ce => 'H',
            sr => \N__50318\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__27869\,
            in2 => \_gnd_net_\,
            in3 => \N__27855\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32111\,
            in1 => \N__28172\,
            in2 => \_gnd_net_\,
            in3 => \N__28158\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__28154\,
            in2 => \_gnd_net_\,
            in3 => \N__28140\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32112\,
            in1 => \N__28136\,
            in2 => \_gnd_net_\,
            in3 => \N__28122\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32085\,
            in1 => \N__28118\,
            in2 => \_gnd_net_\,
            in3 => \N__28104\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32113\,
            in1 => \N__28100\,
            in2 => \_gnd_net_\,
            in3 => \N__28086\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32086\,
            in1 => \N__28082\,
            in2 => \_gnd_net_\,
            in3 => \N__28068\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__28052\,
            in2 => \_gnd_net_\,
            in3 => \N__28038\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__50790\,
            ce => 'H',
            sr => \N__50326\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32115\,
            in1 => \N__28028\,
            in2 => \_gnd_net_\,
            in3 => \N__28014\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32144\,
            in1 => \N__31505\,
            in2 => \_gnd_net_\,
            in3 => \N__28356\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32116\,
            in1 => \N__31529\,
            in2 => \_gnd_net_\,
            in3 => \N__28353\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32145\,
            in1 => \N__28340\,
            in2 => \_gnd_net_\,
            in3 => \N__28326\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32117\,
            in1 => \N__28316\,
            in2 => \_gnd_net_\,
            in3 => \N__28302\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32146\,
            in1 => \N__28289\,
            in2 => \_gnd_net_\,
            in3 => \N__28275\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32118\,
            in1 => \N__28265\,
            in2 => \_gnd_net_\,
            in3 => \N__28251\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32147\,
            in1 => \N__28235\,
            in2 => \_gnd_net_\,
            in3 => \N__28221\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__50781\,
            ce => 'H',
            sr => \N__50334\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32140\,
            in1 => \N__28211\,
            in2 => \_gnd_net_\,
            in3 => \N__28197\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32148\,
            in1 => \N__28192\,
            in2 => \_gnd_net_\,
            in3 => \N__28176\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32141\,
            in1 => \N__28487\,
            in2 => \_gnd_net_\,
            in3 => \N__28473\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32149\,
            in1 => \N__28463\,
            in2 => \_gnd_net_\,
            in3 => \N__28449\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__28439\,
            in2 => \_gnd_net_\,
            in3 => \N__28425\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32150\,
            in1 => \N__28417\,
            in2 => \_gnd_net_\,
            in3 => \N__28398\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32143\,
            in1 => \N__28384\,
            in2 => \_gnd_net_\,
            in3 => \N__28395\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50775\,
            ce => 'H',
            sr => \N__50343\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28681\,
            in2 => \N__31838\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49666\,
            in2 => \N__29745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28362\,
            in2 => \N__49769\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49670\,
            in2 => \N__32952\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32901\,
            in2 => \N__49770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49674\,
            in2 => \N__28536\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28524\,
            in2 => \N__49771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49678\,
            in2 => \N__38544\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49691\,
            in2 => \N__28518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31884\,
            in2 => \N__49775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49679\,
            in2 => \N__28509\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37995\,
            in2 => \N__49772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49683\,
            in2 => \N__30381\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28557\,
            in2 => \N__49773\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49687\,
            in2 => \N__28551\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38319\,
            in2 => \N__49774\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28542\,
            in2 => \N__49776\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49698\,
            in2 => \N__37908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30507\,
            in2 => \N__49777\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49702\,
            in2 => \N__33114\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33258\,
            in2 => \N__49778\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49706\,
            in2 => \N__33060\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28578\,
            in2 => \N__49779\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49710\,
            in2 => \N__30342\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28572\,
            in2 => \N__49780\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49714\,
            in2 => \N__30552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30870\,
            in2 => \N__49781\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49718\,
            in2 => \N__28566\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31083\,
            in2 => \N__49782\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49722\,
            in2 => \N__30753\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29730\,
            in2 => \N__49783\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34340\,
            in2 => \_gnd_net_\,
            in3 => \N__28707\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42836\,
            in1 => \N__42977\,
            in2 => \N__46839\,
            in3 => \N__42236\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28701\,
            in1 => \N__38133\,
            in2 => \N__28704\,
            in3 => \N__31323\,
            lcout => \current_shift_inst.PI_CTRL.N_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42905\,
            in1 => \N__46235\,
            in2 => \N__43865\,
            in3 => \N__42308\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__28695\,
            in1 => \N__34337\,
            in2 => \N__33986\,
            in3 => \N__30605\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31289\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31269\,
            ce => 'H',
            sr => \N__50382\
        );

    \phase_controller_inst2.S2_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50751\,
            ce => \N__43676\,
            sr => \N__50392\
        );

    \phase_controller_inst2.stoper_hc.m10_1_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__34859\,
            in1 => \N__37387\,
            in2 => \_gnd_net_\,
            in3 => \N__31470\,
            lcout => \phase_controller_inst2.stoper_hc.m10Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.m3_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__44126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31469\,
            lcout => \phase_controller_inst2.m3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__37388\,
            in1 => \N__41862\,
            in2 => \N__34812\,
            in3 => \N__34863\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50871\,
            ce => \N__43628\,
            sr => \N__50248\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__29954\,
            in1 => \N__28992\,
            in2 => \_gnd_net_\,
            in3 => \N__29012\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50859\,
            ce => 'H',
            sr => \N__50253\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29120\,
            in1 => \N__29585\,
            in2 => \N__29613\,
            in3 => \N__29102\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28877\,
            in1 => \N__32692\,
            in2 => \_gnd_net_\,
            in3 => \N__28851\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50848\,
            ce => \N__31693\,
            sr => \N__50263\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28802\,
            in1 => \N__32691\,
            in2 => \_gnd_net_\,
            in3 => \N__28779\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50848\,
            ce => \N__31693\,
            sr => \N__50263\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__31427\,
            in1 => \N__29373\,
            in2 => \N__29400\,
            in3 => \N__31418\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__29372\,
            in1 => \N__31428\,
            in2 => \N__31419\,
            in3 => \N__29399\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__29036\,
            in1 => \N__29537\,
            in2 => \N__29052\,
            in3 => \N__29559\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__29121\,
            in1 => \N__29612\,
            in2 => \N__29586\,
            in3 => \N__29103\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.m3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31221\,
            lcout => \phase_controller_inst1.m3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.m37_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__31471\,
            in1 => \N__44081\,
            in2 => \N__44137\,
            in3 => \N__31439\,
            lcout => \phase_controller_inst2.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__29558\,
            in1 => \N__29048\,
            in2 => \N__29538\,
            in3 => \N__29037\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29013\,
            in2 => \N__28955\,
            in3 => \N__28988\,
            lcout => \phase_controller_inst2.stoper_tr.N_38_i\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29943\,
            in1 => \N__28973\,
            in2 => \_gnd_net_\,
            in3 => \N__28959\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29947\,
            in1 => \N__28940\,
            in2 => \N__28956\,
            in3 => \N__28926\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29944\,
            in1 => \N__28922\,
            in2 => \_gnd_net_\,
            in3 => \N__28908\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__28904\,
            in2 => \_gnd_net_\,
            in3 => \N__28890\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29945\,
            in1 => \N__29273\,
            in2 => \_gnd_net_\,
            in3 => \N__29259\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29949\,
            in1 => \N__29252\,
            in2 => \_gnd_net_\,
            in3 => \N__29238\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29946\,
            in1 => \N__29231\,
            in2 => \_gnd_net_\,
            in3 => \N__29217\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__50825\,
            ce => 'H',
            sr => \N__50276\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29953\,
            in1 => \N__29213\,
            in2 => \_gnd_net_\,
            in3 => \N__29199\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29980\,
            in1 => \N__29195\,
            in2 => \_gnd_net_\,
            in3 => \N__29181\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29950\,
            in1 => \N__29177\,
            in2 => \_gnd_net_\,
            in3 => \N__29163\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29981\,
            in1 => \N__29159\,
            in2 => \_gnd_net_\,
            in3 => \N__29145\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29951\,
            in1 => \N__29138\,
            in2 => \_gnd_net_\,
            in3 => \N__29124\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29982\,
            in1 => \N__29444\,
            in2 => \_gnd_net_\,
            in3 => \N__29430\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29952\,
            in1 => \N__29423\,
            in2 => \_gnd_net_\,
            in3 => \N__29409\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29983\,
            in1 => \N__31598\,
            in2 => \_gnd_net_\,
            in3 => \N__29406\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__50815\,
            ce => 'H',
            sr => \N__50286\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29984\,
            in1 => \N__31616\,
            in2 => \_gnd_net_\,
            in3 => \N__29403\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29988\,
            in1 => \N__29390\,
            in2 => \_gnd_net_\,
            in3 => \N__29376\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29985\,
            in1 => \N__29371\,
            in2 => \_gnd_net_\,
            in3 => \N__29355\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29989\,
            in1 => \N__29345\,
            in2 => \_gnd_net_\,
            in3 => \N__29331\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29986\,
            in1 => \N__29318\,
            in2 => \_gnd_net_\,
            in3 => \N__29304\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29990\,
            in1 => \N__29294\,
            in2 => \_gnd_net_\,
            in3 => \N__29280\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29987\,
            in1 => \N__29630\,
            in2 => \_gnd_net_\,
            in3 => \N__29616\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29991\,
            in1 => \N__29608\,
            in2 => \_gnd_net_\,
            in3 => \N__29589\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__50806\,
            ce => 'H',
            sr => \N__50295\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29955\,
            in1 => \N__29581\,
            in2 => \_gnd_net_\,
            in3 => \N__29562\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29959\,
            in1 => \N__29557\,
            in2 => \_gnd_net_\,
            in3 => \N__29541\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29956\,
            in1 => \N__29528\,
            in2 => \_gnd_net_\,
            in3 => \N__29514\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29960\,
            in1 => \N__29509\,
            in2 => \_gnd_net_\,
            in3 => \N__29493\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29957\,
            in1 => \N__29485\,
            in2 => \_gnd_net_\,
            in3 => \N__29469\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29961\,
            in1 => \N__29464\,
            in2 => \_gnd_net_\,
            in3 => \N__29448\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29958\,
            in1 => \N__29837\,
            in2 => \_gnd_net_\,
            in3 => \N__29850\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50798\,
            ce => 'H',
            sr => \N__50302\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39783\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50789\,
            ce => \N__36197\,
            sr => \N__50310\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29760\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__29702\,
            in1 => \N__34330\,
            in2 => \N__29768\,
            in3 => \N__29823\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__38432\,
            in1 => \N__29701\,
            in2 => \_gnd_net_\,
            in3 => \N__29761\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34331\,
            in2 => \_gnd_net_\,
            in3 => \N__30598\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29718\,
            in2 => \N__31865\,
            in3 => \N__31861\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33033\,
            in3 => \N__29649\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32937\,
            in2 => \_gnd_net_\,
            in3 => \N__29646\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32883\,
            in3 => \N__30141\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32889\,
            in2 => \_gnd_net_\,
            in3 => \N__30105\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33045\,
            in2 => \_gnd_net_\,
            in3 => \N__30072\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34947\,
            in2 => \_gnd_net_\,
            in3 => \N__30069\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32847\,
            in2 => \_gnd_net_\,
            in3 => \N__30033\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33039\,
            in2 => \_gnd_net_\,
            in3 => \N__30030\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33156\,
            in2 => \_gnd_net_\,
            in3 => \N__29997\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33195\,
            in2 => \_gnd_net_\,
            in3 => \N__29994\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33099\,
            in2 => \_gnd_net_\,
            in3 => \N__30252\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33093\,
            in2 => \_gnd_net_\,
            in3 => \N__30222\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38073\,
            in2 => \_gnd_net_\,
            in3 => \N__30189\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38121\,
            in2 => \_gnd_net_\,
            in3 => \N__30186\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33024\,
            in2 => \_gnd_net_\,
            in3 => \N__30156\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33183\,
            in3 => \N__30153\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33162\,
            in2 => \_gnd_net_\,
            in3 => \N__30150\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33168\,
            in2 => \_gnd_net_\,
            in3 => \N__30147\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33150\,
            in2 => \_gnd_net_\,
            in3 => \N__30144\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33174\,
            in2 => \_gnd_net_\,
            in3 => \N__30333\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33246\,
            in2 => \_gnd_net_\,
            in3 => \N__30303\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33303\,
            in2 => \_gnd_net_\,
            in3 => \N__30300\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33189\,
            in2 => \_gnd_net_\,
            in3 => \N__30297\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33297\,
            in2 => \_gnd_net_\,
            in3 => \N__30294\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33144\,
            in2 => \_gnd_net_\,
            in3 => \N__30291\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33291\,
            in2 => \_gnd_net_\,
            in3 => \N__30261\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36090\,
            in2 => \_gnd_net_\,
            in3 => \N__30258\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__30255\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30615\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34225\,
            in1 => \N__35641\,
            in2 => \_gnd_net_\,
            in3 => \N__30568\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38524\,
            in1 => \N__35386\,
            in2 => \_gnd_net_\,
            in3 => \N__30523\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__30498\,
            in1 => \N__30486\,
            in2 => \_gnd_net_\,
            in3 => \N__34726\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34727\,
            in1 => \N__30477\,
            in2 => \_gnd_net_\,
            in3 => \N__30468\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__30456\,
            in1 => \N__30444\,
            in2 => \_gnd_net_\,
            in3 => \N__34728\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__34729\,
            in1 => \N__30435\,
            in2 => \_gnd_net_\,
            in3 => \N__30423\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38522\,
            in1 => \N__35527\,
            in2 => \_gnd_net_\,
            in3 => \N__30406\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35737\,
            in1 => \N__38523\,
            in2 => \_gnd_net_\,
            in3 => \N__30364\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__30816\,
            in1 => \N__30804\,
            in2 => \_gnd_net_\,
            in3 => \N__34730\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__36067\,
            in1 => \N__34314\,
            in2 => \_gnd_net_\,
            in3 => \N__30769\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34699\,
            in1 => \N__30741\,
            in2 => \_gnd_net_\,
            in3 => \N__30732\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__30720\,
            in1 => \N__30711\,
            in2 => \_gnd_net_\,
            in3 => \N__34697\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30699\,
            in3 => \N__33233\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50765\,
            ce => 'H',
            sr => \N__50355\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34698\,
            lcout => \current_shift_inst.N_1275_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34700\,
            in1 => \N__30660\,
            in2 => \_gnd_net_\,
            in3 => \N__30648\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__30636\,
            in1 => \N__30627\,
            in2 => \_gnd_net_\,
            in3 => \N__34701\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34708\,
            in1 => \N__31047\,
            in2 => \_gnd_net_\,
            in3 => \N__31035\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__31023\,
            in1 => \N__31011\,
            in2 => \_gnd_net_\,
            in3 => \N__34709\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__34710\,
            in1 => \_gnd_net_\,
            in2 => \N__30999\,
            in3 => \N__30984\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__30969\,
            in1 => \N__30960\,
            in2 => \_gnd_net_\,
            in3 => \N__34711\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__34712\,
            in1 => \N__30948\,
            in2 => \_gnd_net_\,
            in3 => \N__30936\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__30924\,
            in1 => \N__30912\,
            in2 => \_gnd_net_\,
            in3 => \N__34707\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34312\,
            in1 => \N__35602\,
            in2 => \_gnd_net_\,
            in3 => \N__30889\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__30861\,
            in1 => \N__30849\,
            in2 => \_gnd_net_\,
            in3 => \N__34706\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__30840\,
            in1 => \N__30828\,
            in2 => \_gnd_net_\,
            in3 => \N__34719\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__34720\,
            in1 => \N__31182\,
            in2 => \_gnd_net_\,
            in3 => \N__31170\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31158\,
            in1 => \N__31146\,
            in2 => \_gnd_net_\,
            in3 => \N__34718\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__34721\,
            in1 => \N__31134\,
            in2 => \_gnd_net_\,
            in3 => \N__31122\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__36121\,
            in1 => \N__34313\,
            in2 => \_gnd_net_\,
            in3 => \N__31108\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34722\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31071\,
            in1 => \N__31062\,
            in2 => \_gnd_net_\,
            in3 => \N__34740\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43514\,
            in1 => \N__42719\,
            in2 => \N__43358\,
            in3 => \N__42772\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43915\,
            in1 => \N__43978\,
            in2 => \N__43802\,
            in3 => \N__43165\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__43231\,
            in1 => \N__43466\,
            in2 => \N__31050\,
            in3 => \N__31317\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__43282\,
            in1 => \N__46585\,
            in2 => \N__31332\,
            in3 => \N__31329\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43106\,
            in2 => \_gnd_net_\,
            in3 => \N__43402\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31288\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__31268\,
            ce => 'H',
            sr => \N__50378\
        );

    \phase_controller_inst2.S1_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41918\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50750\,
            ce => \N__43663\,
            sr => \N__50387\
        );

    \GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_red_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_0_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__37463\,
            in1 => \N__37533\,
            in2 => \N__38845\,
            in3 => \N__40642\,
            lcout => \phase_controller_inst1.stoper_hc.m19_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_1_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__37534\,
            in2 => \N__38856\,
            in3 => \N__40635\,
            lcout => \phase_controller_inst1.stoper_hc.m34_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__37584\,
            in1 => \N__34933\,
            in2 => \N__31213\,
            in3 => \N__31230\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50882\,
            ce => \N__43627\,
            sr => \N__50244\
        );

    \phase_controller_inst2.start_timer_tr_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__42152\,
            in1 => \N__34906\,
            in2 => \N__44208\,
            in3 => \N__31188\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50882\,
            ce => \N__43627\,
            sr => \N__50244\
        );

    \phase_controller_inst2.state_1_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__34878\,
            in1 => \N__34864\,
            in2 => \N__37401\,
            in3 => \N__34907\,
            lcout => \phase_controller_inst2.N_139_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50882\,
            ce => \N__43627\,
            sr => \N__50244\
        );

    \phase_controller_inst2.stoper_hc.m20_ns_1_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001000"
        )
    port map (
            in0 => \N__42115\,
            in1 => \N__41908\,
            in2 => \N__44204\,
            in3 => \N__34904\,
            lcout => \phase_controller_inst2.stoper_hc.m20_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__34995\,
            in1 => \N__48171\,
            in2 => \N__51520\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50861\,
            ce => \N__49248\,
            sr => \N__50254\
        );

    \phase_controller_inst2.stoper_hc.m38_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101110101"
        )
    port map (
            in0 => \N__31472\,
            in1 => \N__44082\,
            in2 => \N__44144\,
            in3 => \N__31443\,
            lcout => \phase_controller_inst2.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32669\,
            in1 => \N__32252\,
            in2 => \_gnd_net_\,
            in3 => \N__32232\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32767\,
            in1 => \N__32748\,
            in2 => \_gnd_net_\,
            in3 => \N__32668\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32248\,
            in1 => \N__32231\,
            in2 => \_gnd_net_\,
            in3 => \N__32563\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50840\,
            ce => \N__31699\,
            sr => \N__50270\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32821\,
            in1 => \N__32562\,
            in2 => \_gnd_net_\,
            in3 => \N__32841\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50840\,
            ce => \N__31699\,
            sr => \N__50270\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__31407\,
            in2 => \_gnd_net_\,
            in3 => \N__31365\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50827\,
            ce => \N__31701\,
            sr => \N__50277\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31815\,
            in1 => \N__31782\,
            in2 => \_gnd_net_\,
            in3 => \N__32690\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50827\,
            ce => \N__31701\,
            sr => \N__50277\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32688\,
            in1 => \N__31767\,
            in2 => \_gnd_net_\,
            in3 => \N__31746\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50827\,
            ce => \N__31701\,
            sr => \N__50277\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__41300\,
            in1 => \N__41552\,
            in2 => \N__31650\,
            in3 => \N__31662\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__31661\,
            in1 => \N__41301\,
            in2 => \N__41553\,
            in3 => \N__31646\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34973\,
            in1 => \_gnd_net_\,
            in2 => \N__51516\,
            in3 => \N__45057\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50817\,
            ce => \N__49241\,
            sr => \N__50287\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__31594\,
            in1 => \N__31578\,
            in2 => \N__31617\,
            in3 => \N__31626\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__31625\,
            in1 => \N__31615\,
            in2 => \N__31599\,
            in3 => \N__31577\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__31536\,
            in1 => \N__31511\,
            in2 => \N__32784\,
            in3 => \N__32187\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__32186\,
            in1 => \N__31535\,
            in2 => \N__31515\,
            in3 => \N__32780\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32822\,
            in1 => \N__32684\,
            in2 => \_gnd_net_\,
            in3 => \N__32837\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32686\,
            in1 => \_gnd_net_\,
            in2 => \N__32826\,
            in3 => \N__32823\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50808\,
            ce => \N__32139\,
            sr => \N__50296\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32772\,
            in1 => \N__32746\,
            in2 => \_gnd_net_\,
            in3 => \N__32687\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50808\,
            ce => \N__32139\,
            sr => \N__50296\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32685\,
            in1 => \N__32253\,
            in2 => \_gnd_net_\,
            in3 => \N__32230\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50808\,
            ce => \N__32139\,
            sr => \N__50296\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34332\,
            in2 => \_gnd_net_\,
            in3 => \N__33975\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35086\,
            in1 => \N__38431\,
            in2 => \_gnd_net_\,
            in3 => \N__31909\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33001\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__33002\,
            in1 => \_gnd_net_\,
            in2 => \N__31842\,
            in3 => \N__38430\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36160\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50800\,
            ce => \N__36195\,
            sr => \N__50303\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39456\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50800\,
            ce => \N__36195\,
            sr => \N__50303\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35296\,
            in1 => \N__38447\,
            in2 => \_gnd_net_\,
            in3 => \N__32968\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35295\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__38448\,
            in2 => \_gnd_net_\,
            in3 => \N__32917\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35210\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35259\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32874\,
            in1 => \N__32862\,
            in2 => \_gnd_net_\,
            in3 => \N__34752\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35113\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38497\,
            in1 => \N__35917\,
            in2 => \_gnd_net_\,
            in3 => \N__33130\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35508\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35464\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.m16_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34911\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42132\,
            lcout => \phase_controller_inst2.stoper_hc.mZ0Z16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38498\,
            in1 => \N__35833\,
            in2 => \_gnd_net_\,
            in3 => \N__33076\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35164\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35072\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35327\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35413\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38047\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37960\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35823\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35376\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35035\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35863\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35588\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__34311\,
            in1 => \N__35683\,
            in2 => \N__33990\,
            in3 => \N__33343\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35718\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35555\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35864\,
            in1 => \N__38525\,
            in2 => \_gnd_net_\,
            in3 => \N__33269\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35767\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33240\,
            in2 => \N__33234\,
            in3 => \N__33232\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33213\,
            in2 => \_gnd_net_\,
            in3 => \N__33207\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33204\,
            in2 => \_gnd_net_\,
            in3 => \N__33198\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34425\,
            in2 => \_gnd_net_\,
            in3 => \N__34419\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34416\,
            in2 => \_gnd_net_\,
            in3 => \N__34410\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34407\,
            in2 => \_gnd_net_\,
            in3 => \N__34395\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34392\,
            in2 => \_gnd_net_\,
            in3 => \N__34386\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34383\,
            in2 => \_gnd_net_\,
            in3 => \N__34371\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34368\,
            in2 => \_gnd_net_\,
            in3 => \N__34362\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34359\,
            in2 => \_gnd_net_\,
            in3 => \N__34353\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34350\,
            in2 => \_gnd_net_\,
            in3 => \N__34344\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34506\,
            in2 => \_gnd_net_\,
            in3 => \N__34500\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34497\,
            in2 => \_gnd_net_\,
            in3 => \N__34491\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34488\,
            in2 => \_gnd_net_\,
            in3 => \N__34482\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34479\,
            in2 => \_gnd_net_\,
            in3 => \N__34473\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34470\,
            in2 => \_gnd_net_\,
            in3 => \N__34464\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34461\,
            in2 => \_gnd_net_\,
            in3 => \N__34452\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34449\,
            in2 => \_gnd_net_\,
            in3 => \N__34443\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34440\,
            in3 => \N__34428\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34599\,
            in2 => \_gnd_net_\,
            in3 => \N__34590\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34587\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34578\,
            in2 => \_gnd_net_\,
            in3 => \N__34572\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34569\,
            in2 => \_gnd_net_\,
            in3 => \N__34563\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34560\,
            in2 => \_gnd_net_\,
            in3 => \N__34554\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34551\,
            in2 => \_gnd_net_\,
            in3 => \N__34542\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34539\,
            in2 => \_gnd_net_\,
            in3 => \N__34533\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34530\,
            in2 => \_gnd_net_\,
            in3 => \N__34521\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34518\,
            in2 => \_gnd_net_\,
            in3 => \N__34509\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34773\,
            in2 => \_gnd_net_\,
            in3 => \N__34764\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34761\,
            in2 => \_gnd_net_\,
            in3 => \N__34755\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34751\,
            in2 => \_gnd_net_\,
            in3 => \N__34602\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42018\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50758\,
            ce => 'H',
            sr => \N__50365\
        );

    \phase_controller_inst2.stoper_hc.running_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__42045\,
            in1 => \N__42083\,
            in2 => \_gnd_net_\,
            in3 => \N__41984\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50758\,
            ce => 'H',
            sr => \N__50365\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37115\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__46589\,
            in1 => \N__46378\,
            in2 => \N__42402\,
            in3 => \N__46780\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50757\,
            ce => 'H',
            sr => \N__50372\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__42017\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42049\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_RNI3USR_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__34937\,
            in1 => \N__38832\,
            in2 => \N__40643\,
            in3 => \N__37575\,
            lcout => \phase_controller_inst1.stoper_hc.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_RNI61TR_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000110001001"
        )
    port map (
            in0 => \N__38820\,
            in1 => \N__38773\,
            in2 => \N__34938\,
            in3 => \N__40631\,
            lcout => \phase_controller_inst1.stoper_hc.m12_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_er_RNI72V01_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__34808\,
            in1 => \N__44203\,
            in2 => \N__41858\,
            in3 => \N__34905\,
            lcout => \phase_controller_inst2.stoper_hc.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.m21_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41892\,
            lcout => \phase_controller_inst2.m21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_er_RNI23UO1_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001001111"
        )
    port map (
            in0 => \N__34804\,
            in1 => \N__41891\,
            in2 => \N__41857\,
            in3 => \N__34872\,
            lcout => \phase_controller_inst2.time_passed_er_RNI23UO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_er_RNI0D511_0_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111010011"
        )
    port map (
            in0 => \N__34803\,
            in1 => \N__37402\,
            in2 => \N__41856\,
            in3 => \N__34866\,
            lcout => \phase_controller_inst2.stoper_hc.m28_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_er_RNI7HLK_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34799\,
            in2 => \_gnd_net_\,
            in3 => \N__41843\,
            lcout => \phase_controller_inst2.stoper_hc.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_er_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42069\,
            lcout => \phase_controller_inst2.stoper_hc.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50862\,
            ce => \N__35004\,
            sr => \N__50255\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__35016\,
            in1 => \N__37697\,
            in2 => \N__37830\,
            in3 => \N__37720\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39535\,
            in1 => \N__44679\,
            in2 => \_gnd_net_\,
            in3 => \N__51299\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50850\,
            ce => \N__48826\,
            sr => \N__50264\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51285\,
            in1 => \N__34974\,
            in2 => \_gnd_net_\,
            in3 => \N__45055\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101110001"
        )
    port map (
            in0 => \N__37722\,
            in1 => \N__37696\,
            in2 => \N__37826\,
            in3 => \N__35015\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51284\,
            in1 => \N__48163\,
            in2 => \_gnd_net_\,
            in3 => \N__34994\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_sbtinv_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41988\,
            lcout => \phase_controller_inst2.stoper_hc.N_266_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44678\,
            in1 => \N__39539\,
            in2 => \_gnd_net_\,
            in3 => \N__51283\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34990\,
            in1 => \N__48170\,
            in2 => \_gnd_net_\,
            in3 => \N__51300\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50828\,
            ce => \N__48862\,
            sr => \N__50278\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34972\,
            in1 => \N__45056\,
            in2 => \_gnd_net_\,
            in3 => \N__51301\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50828\,
            ce => \N__48862\,
            sr => \N__50278\
        );

    \delay_measurement_inst.start_timer_hc_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34956\,
            ce => 'H',
            sr => \N__50288\
        );

    \delay_measurement_inst.stop_timer_hc_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38271\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34956\,
            ce => 'H',
            sr => \N__50288\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38592\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39749\,
            in2 => \N__39455\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39728\,
            in2 => \N__39782\,
            in3 => \N__35277\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39750\,
            in2 => \N__39707\,
            in3 => \N__35241\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39729\,
            in2 => \N__39680\,
            in3 => \N__35199\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39653\,
            in2 => \N__39708\,
            in3 => \N__35148\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39632\,
            in2 => \N__39681\,
            in3 => \N__35145\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39654\,
            in2 => \N__39611\,
            in3 => \N__35097\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39633\,
            in2 => \N__40026\,
            in3 => \N__35061\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__50791\,
            ce => \N__36194\,
            sr => \N__50311\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39989\,
            in2 => \N__39612\,
            in3 => \N__35019\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39968\,
            in2 => \N__40025\,
            in3 => \N__35541\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39990\,
            in2 => \N__39948\,
            in3 => \N__35490\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39969\,
            in2 => \N__39920\,
            in3 => \N__35448\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39947\,
            in2 => \N__39893\,
            in3 => \N__35445\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39866\,
            in2 => \N__39921\,
            in3 => \N__35442\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39842\,
            in2 => \N__39894\,
            in3 => \N__35400\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39867\,
            in2 => \N__39815\,
            in3 => \N__35397\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__50782\,
            ce => \N__36193\,
            sr => \N__50319\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40238\,
            in2 => \N__39846\,
            in3 => \N__35358\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40217\,
            in2 => \N__39816\,
            in3 => \N__35889\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40239\,
            in2 => \N__40194\,
            in3 => \N__35847\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40218\,
            in2 => \N__40167\,
            in3 => \N__35805\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40193\,
            in2 => \N__40139\,
            in3 => \N__35751\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40166\,
            in2 => \N__40112\,
            in3 => \N__35697\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40082\,
            in2 => \N__40140\,
            in3 => \N__35661\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40052\,
            in2 => \N__40113\,
            in3 => \N__35616\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__50776\,
            ce => \N__36192\,
            sr => \N__50327\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40406\,
            in2 => \N__40086\,
            in3 => \N__35577\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__50771\,
            ce => \N__36191\,
            sr => \N__50335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40382\,
            in2 => \N__40056\,
            in3 => \N__35544\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__50771\,
            ce => \N__36191\,
            sr => \N__50335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40362\,
            in2 => \N__40410\,
            in3 => \N__36204\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__50771\,
            ce => \N__36191\,
            sr => \N__50335\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40383\,
            in2 => \N__40341\,
            in3 => \N__36201\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__50771\,
            ce => \N__36191\,
            sr => \N__50335\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36168\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36103\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36058\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36027\,
            in2 => \_gnd_net_\,
            in3 => \N__36033\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36021\,
            in2 => \_gnd_net_\,
            in3 => \N__35979\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35976\,
            in2 => \_gnd_net_\,
            in3 => \N__35940\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36456\,
            in2 => \_gnd_net_\,
            in3 => \N__36417\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36414\,
            in2 => \_gnd_net_\,
            in3 => \N__36408\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36405\,
            in2 => \_gnd_net_\,
            in3 => \N__36372\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36369\,
            in2 => \_gnd_net_\,
            in3 => \N__36330\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36327\,
            in2 => \_gnd_net_\,
            in3 => \N__36300\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__50770\,
            ce => 'H',
            sr => \N__50344\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36297\,
            in2 => \_gnd_net_\,
            in3 => \N__36291\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36288\,
            in2 => \_gnd_net_\,
            in3 => \N__36249\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36246\,
            in2 => \_gnd_net_\,
            in3 => \N__36207\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36774\,
            in2 => \_gnd_net_\,
            in3 => \N__36735\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36732\,
            in2 => \_gnd_net_\,
            in3 => \N__36693\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36690\,
            in2 => \_gnd_net_\,
            in3 => \N__36657\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36654\,
            in2 => \_gnd_net_\,
            in3 => \N__36621\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36618\,
            in2 => \_gnd_net_\,
            in3 => \N__36588\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__50768\,
            ce => 'H',
            sr => \N__50350\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36585\,
            in2 => \_gnd_net_\,
            in3 => \N__36540\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36537\,
            in2 => \_gnd_net_\,
            in3 => \N__36504\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36501\,
            in2 => \_gnd_net_\,
            in3 => \N__36459\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37065\,
            in2 => \_gnd_net_\,
            in3 => \N__37032\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37029\,
            in2 => \_gnd_net_\,
            in3 => \N__36993\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36990\,
            in2 => \_gnd_net_\,
            in3 => \N__36951\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36948\,
            in2 => \_gnd_net_\,
            in3 => \N__36915\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36912\,
            in2 => \_gnd_net_\,
            in3 => \N__36879\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__50766\,
            ce => 'H',
            sr => \N__50356\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36876\,
            in2 => \_gnd_net_\,
            in3 => \N__36831\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36828\,
            in2 => \_gnd_net_\,
            in3 => \N__36783\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36780\,
            in2 => \_gnd_net_\,
            in3 => \N__37284\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37281\,
            in2 => \_gnd_net_\,
            in3 => \N__37239\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37236\,
            in2 => \_gnd_net_\,
            in3 => \N__37197\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37194\,
            in2 => \_gnd_net_\,
            in3 => \N__37158\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37155\,
            in2 => \_gnd_net_\,
            in3 => \N__37119\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37116\,
            in2 => \_gnd_net_\,
            in3 => \N__37104\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50762\,
            ce => 'H',
            sr => \N__50361\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__46750\,
            in1 => \N__46597\,
            in2 => \N__42600\,
            in3 => \N__46379\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50759\,
            ce => 'H',
            sr => \N__50366\
        );

    \phase_controller_inst1.S2_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37479\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50756\,
            ce => \N__43659\,
            sr => \N__50379\
        );

    \phase_controller_inst1.state_3_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__38787\,
            in1 => \N__37580\,
            in2 => \N__38855\,
            in3 => \N__37074\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50907\,
            ce => \N__43599\,
            sr => \N__50229\
        );

    \phase_controller_inst1.state_1_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__37541\,
            in1 => \N__37579\,
            in2 => \N__37471\,
            in3 => \N__37605\,
            lcout => \phase_controller_inst1.N_175_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50907\,
            ce => \N__43599\,
            sr => \N__50229\
        );

    \phase_controller_inst1.state_2_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110100000"
        )
    port map (
            in0 => \N__38833\,
            in1 => \N__37542\,
            in2 => \N__40644\,
            in3 => \N__37462\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50907\,
            ce => \N__43599\,
            sr => \N__50229\
        );

    \phase_controller_inst1.stoper_hc.m7_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37599\,
            in2 => \_gnd_net_\,
            in3 => \N__38770\,
            lcout => \phase_controller_inst1.stoper_hc.N_8_0\,
            ltout => \phase_controller_inst1.stoper_hc.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_RNINITI1_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100100011"
        )
    port map (
            in0 => \N__37574\,
            in1 => \N__38844\,
            in2 => \N__37551\,
            in3 => \N__37548\,
            lcout => \phase_controller_inst1.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.m13_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__38772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37540\,
            lcout => \phase_controller_inst1.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_RNI9RLH_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__38771\,
            in1 => \N__43626\,
            in2 => \_gnd_net_\,
            in3 => \N__37328\,
            lcout => \S1_RNI9RLH\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__37497\,
            in1 => \N__38702\,
            in2 => \N__37491\,
            in3 => \N__37470\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50897\,
            ce => \N__43607\,
            sr => \N__50237\
        );

    \phase_controller_inst2.state_4_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__38714\,
            in1 => \N__37422\,
            in2 => \N__37415\,
            in3 => \N__37353\,
            lcout => \phase_controller_inst2.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50897\,
            ce => \N__43607\,
            sr => \N__50237\
        );

    \phase_controller_inst1.S1_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38775\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50897\,
            ce => \N__43607\,
            sr => \N__50237\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40575\,
            in2 => \N__37640\,
            in3 => \N__40586\,
            lcout => \phase_controller_inst1.stoper_hc.N_45_i\,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48712\,
            in1 => \N__39024\,
            in2 => \_gnd_net_\,
            in3 => \N__37644\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__48809\,
            in1 => \N__39003\,
            in2 => \N__37641\,
            in3 => \N__37626\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48713\,
            in1 => \N__38985\,
            in2 => \_gnd_net_\,
            in3 => \N__37623\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48810\,
            in1 => \N__38964\,
            in2 => \_gnd_net_\,
            in3 => \N__37620\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48714\,
            in1 => \N__38931\,
            in2 => \_gnd_net_\,
            in3 => \N__37617\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48811\,
            in1 => \N__38898\,
            in2 => \_gnd_net_\,
            in3 => \N__37614\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48715\,
            in1 => \N__38877\,
            in2 => \_gnd_net_\,
            in3 => \N__37611\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50890\,
            ce => 'H',
            sr => \N__50240\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48723\,
            in1 => \N__39189\,
            in2 => \_gnd_net_\,
            in3 => \N__37608\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48716\,
            in1 => \N__39171\,
            in2 => \_gnd_net_\,
            in3 => \N__37671\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48720\,
            in1 => \N__39150\,
            in2 => \_gnd_net_\,
            in3 => \N__37668\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48717\,
            in1 => \N__39129\,
            in2 => \_gnd_net_\,
            in3 => \N__37665\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48721\,
            in1 => \N__39102\,
            in2 => \_gnd_net_\,
            in3 => \N__37662\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48718\,
            in1 => \N__39078\,
            in2 => \_gnd_net_\,
            in3 => \N__37659\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48722\,
            in1 => \N__39045\,
            in2 => \_gnd_net_\,
            in3 => \N__37656\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48719\,
            in1 => \N__40795\,
            in2 => \_gnd_net_\,
            in3 => \N__37653\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__50883\,
            ce => 'H',
            sr => \N__50245\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48838\,
            in1 => \N__40811\,
            in2 => \_gnd_net_\,
            in3 => \N__37650\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48751\,
            in1 => \N__39331\,
            in2 => \_gnd_net_\,
            in3 => \N__37647\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48839\,
            in1 => \N__39352\,
            in2 => \_gnd_net_\,
            in3 => \N__37737\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48752\,
            in1 => \N__39389\,
            in2 => \_gnd_net_\,
            in3 => \N__37734\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48840\,
            in1 => \N__39412\,
            in2 => \_gnd_net_\,
            in3 => \N__37731\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48753\,
            in1 => \N__40859\,
            in2 => \_gnd_net_\,
            in3 => \N__37728\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48841\,
            in1 => \N__40880\,
            in2 => \_gnd_net_\,
            in3 => \N__37725\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48754\,
            in1 => \N__37721\,
            in2 => \_gnd_net_\,
            in3 => \N__37701\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__50873\,
            ce => 'H',
            sr => \N__50249\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48842\,
            in1 => \N__37698\,
            in2 => \_gnd_net_\,
            in3 => \N__37680\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48833\,
            in1 => \N__40691\,
            in2 => \_gnd_net_\,
            in3 => \N__37677\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48843\,
            in1 => \N__40670\,
            in2 => \_gnd_net_\,
            in3 => \N__37674\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48834\,
            in1 => \N__37879\,
            in2 => \_gnd_net_\,
            in3 => \N__37803\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48844\,
            in1 => \N__37858\,
            in2 => \_gnd_net_\,
            in3 => \N__37800\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48835\,
            in1 => \N__37791\,
            in2 => \_gnd_net_\,
            in3 => \N__37797\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__37775\,
            in1 => \N__48836\,
            in2 => \_gnd_net_\,
            in3 => \N__37794\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50863\,
            ce => 'H',
            sr => \N__50256\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51386\,
            in1 => \N__49201\,
            in2 => \_gnd_net_\,
            in3 => \N__49164\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50851\,
            ce => \N__48837\,
            sr => \N__50265\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__37745\,
            in1 => \N__37790\,
            in2 => \N__37776\,
            in3 => \N__37754\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__37789\,
            in1 => \N__37774\,
            in2 => \N__37758\,
            in3 => \N__37746\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42187\,
            in1 => \N__44985\,
            in2 => \_gnd_net_\,
            in3 => \N__51387\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50851\,
            ce => \N__48837\,
            sr => \N__50265\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__48126\,
            in1 => \N__49200\,
            in2 => \N__47781\,
            in3 => \N__39285\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44481\,
            in2 => \N__37893\,
            in3 => \N__44349\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50851\,
            ce => \N__48837\,
            sr => \N__50265\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__37880\,
            in1 => \N__37890\,
            in2 => \N__37842\,
            in3 => \N__37862\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__37889\,
            in1 => \N__37881\,
            in2 => \N__37863\,
            in3 => \N__37841\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47853\,
            in1 => \N__39477\,
            in2 => \_gnd_net_\,
            in3 => \N__51298\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50841\,
            ce => \N__48866\,
            sr => \N__50271\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51389\,
            in1 => \N__39517\,
            in2 => \_gnd_net_\,
            in3 => \N__48215\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50829\,
            ce => \N__48851\,
            sr => \N__50279\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45347\,
            in1 => \N__45364\,
            in2 => \_gnd_net_\,
            in3 => \N__51390\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50829\,
            ce => \N__48851\,
            sr => \N__50279\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51388\,
            in1 => \N__39577\,
            in2 => \_gnd_net_\,
            in3 => \N__44618\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50829\,
            ce => \N__48851\,
            sr => \N__50279\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44806\,
            in1 => \N__39559\,
            in2 => \_gnd_net_\,
            in3 => \N__51391\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50829\,
            ce => \N__48851\,
            sr => \N__50279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39561\,
            in1 => \N__44805\,
            in2 => \_gnd_net_\,
            in3 => \N__51318\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38252\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51415\,
            in1 => \N__47855\,
            in2 => \_gnd_net_\,
            in3 => \N__39476\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38253\,
            in2 => \_gnd_net_\,
            in3 => \N__38296\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_341_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38376\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNI419P_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__38178\,
            in1 => \N__49130\,
            in2 => \_gnd_net_\,
            in3 => \N__38679\,
            lcout => \current_shift_inst.timer_s1.N_340_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38084\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38185\,
            in2 => \_gnd_net_\,
            in3 => \N__38153\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50792\,
            ce => 'H',
            sr => \N__50312\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38519\,
            in1 => \N__38048\,
            in2 => \_gnd_net_\,
            in3 => \N__38029\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38520\,
            in1 => \N__37961\,
            in2 => \_gnd_net_\,
            in3 => \N__37933\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38518\,
            in1 => \N__38602\,
            in2 => \_gnd_net_\,
            in3 => \N__38569\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__38279\,
            in1 => \N__38250\,
            in2 => \_gnd_net_\,
            in3 => \N__38303\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_342_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38521\,
            in1 => \N__38377\,
            in2 => \_gnd_net_\,
            in3 => \N__38351\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__38251\,
            in1 => \N__38304\,
            in2 => \_gnd_net_\,
            in3 => \N__38280\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50777\,
            ce => 'H',
            sr => \N__50328\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38222\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50777\,
            ce => 'H',
            sr => \N__50328\
        );

    \current_shift_inst.timer_s1.running_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__38186\,
            in1 => \N__49119\,
            in2 => \_gnd_net_\,
            in3 => \N__38678\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50777\,
            ce => 'H',
            sr => \N__50328\
        );

    \current_shift_inst.stop_timer_s1_er_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38187\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50772\,
            ce => \N__38160\,
            sr => \N__50336\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__41627\,
            in1 => \N__41692\,
            in2 => \N__41794\,
            in3 => \N__42654\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__40248\,
            in1 => \N__42374\,
            in2 => \N__38136\,
            in3 => \N__46891\,
            lcout => \current_shift_inst.PI_CTRL.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNI8ENL_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49120\,
            in2 => \_gnd_net_\,
            in3 => \N__38674\,
            lcout => \current_shift_inst.timer_s1.N_339_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46556\,
            in1 => \N__43403\,
            in2 => \N__43232\,
            in3 => \N__43462\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42893\,
            in1 => \N__46234\,
            in2 => \N__42301\,
            in3 => \N__42835\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46825\,
            in1 => \N__43801\,
            in2 => \N__38640\,
            in3 => \N__38622\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38637\,
            in1 => \N__38628\,
            in2 => \N__38631\,
            in3 => \N__40422\,
            lcout => \current_shift_inst.PI_CTRL.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43979\,
            in1 => \N__43166\,
            in2 => \N__43922\,
            in3 => \N__43096\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42958\,
            in2 => \_gnd_net_\,
            in3 => \N__42226\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__46748\,
            in1 => \N__41777\,
            in2 => \N__41742\,
            in3 => \N__46374\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50763\,
            ce => 'H',
            sr => \N__50362\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__46372\,
            in1 => \N__46545\,
            in2 => \N__42684\,
            in3 => \N__46749\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50763\,
            ce => 'H',
            sr => \N__50362\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__46544\,
            in1 => \N__46373\,
            in2 => \N__46781\,
            in3 => \N__43425\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50763\,
            ce => 'H',
            sr => \N__50362\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__41646\,
            in1 => \N__46418\,
            in2 => \_gnd_net_\,
            in3 => \N__46751\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50760\,
            ce => 'H',
            sr => \N__50367\
        );

    \phase_controller_inst1.start_timer_hc_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__38834\,
            in1 => \N__40615\,
            in2 => \N__40554\,
            in3 => \N__38786\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50908\,
            ce => \N__43625\,
            sr => \N__50230\
        );

    \phase_controller_inst1.test22_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__43606\,
            in1 => \N__38726\,
            in2 => \_gnd_net_\,
            in3 => \N__38774\,
            lcout => test22_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50902\,
            ce => 'H',
            sr => \N__50233\
        );

    \phase_controller_inst2.state_0_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38715\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50902\,
            ce => 'H',
            sr => \N__50233\
        );

    \phase_controller_inst1.state_0_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38703\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50902\,
            ce => 'H',
            sr => \N__50233\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40550\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50902\,
            ce => 'H',
            sr => \N__50233\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_0_30_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__40551\,
            in1 => \N__40511\,
            in2 => \N__40487\,
            in3 => \N__40463\,
            lcout => \phase_controller_inst1.stoper_hc.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__40512\,
            in1 => \N__40552\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44016\,
            in2 => \N__38691\,
            in3 => \N__40570\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47931\,
            in2 => \N__39012\,
            in3 => \N__39023\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38991\,
            in2 => \N__44157\,
            in3 => \N__39002\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40752\,
            in2 => \N__38973\,
            in3 => \N__38984\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40710\,
            in2 => \N__38952\,
            in3 => \N__38963\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38943\,
            in2 => \N__38919\,
            in3 => \N__38930\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38910\,
            in2 => \N__38886\,
            in3 => \N__38897\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44028\,
            in2 => \N__38865\,
            in3 => \N__38876\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39188\,
            in1 => \N__39177\,
            in2 => \N__47919\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40716\,
            in2 => \N__39159\,
            in3 => \N__39170\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47907\,
            in2 => \N__39138\,
            in3 => \N__39149\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39117\,
            in2 => \N__40725\,
            in3 => \N__39128\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39111\,
            in2 => \N__39090\,
            in3 => \N__39101\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39306\,
            in2 => \N__39066\,
            in3 => \N__39077\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39057\,
            in2 => \N__39033\,
            in3 => \N__39044\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40824\,
            in2 => \N__40770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39315\,
            in2 => \N__39198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39375\,
            in2 => \N__39279\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40845\,
            in2 => \N__40908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39267\,
            in2 => \N__39258\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40650\,
            in2 => \N__40704\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39243\,
            in2 => \N__39231\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39216\,
            in2 => \N__39210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39201\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__39354\,
            in1 => \N__47969\,
            in2 => \N__39336\,
            in3 => \N__39297\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__39296\,
            in1 => \N__39353\,
            in2 => \N__47973\,
            in3 => \N__39335\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45425\,
            in1 => \N__45383\,
            in2 => \_gnd_net_\,
            in3 => \N__51280\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51281\,
            in1 => \_gnd_net_\,
            in2 => \N__39309\,
            in3 => \N__45426\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50864\,
            ce => \N__48825\,
            sr => \N__50257\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45275\,
            in1 => \N__45252\,
            in2 => \_gnd_net_\,
            in3 => \N__51282\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50864\,
            ce => \N__48825\,
            sr => \N__50257\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45045\,
            in1 => \N__45183\,
            in2 => \N__44619\,
            in3 => \N__44982\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39360\,
            in1 => \N__39366\,
            in2 => \N__39288\,
            in3 => \N__44004\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42191\,
            in1 => \N__51317\,
            in2 => \_gnd_net_\,
            in3 => \N__44983\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__39423\,
            in1 => \N__39414\,
            in2 => \N__48894\,
            in3 => \N__39396\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51287\,
            in1 => \N__48961\,
            in2 => \_gnd_net_\,
            in3 => \N__48936\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__39422\,
            in1 => \N__39413\,
            in2 => \N__48893\,
            in3 => \N__39395\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51286\,
            in1 => \N__45493\,
            in2 => \_gnd_net_\,
            in3 => \N__45470\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__39518\,
            in1 => \_gnd_net_\,
            in2 => \N__48214\,
            in3 => \N__51288\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51123\,
            in1 => \N__51763\,
            in2 => \N__48939\,
            in3 => \N__44671\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49473\,
            in1 => \N__45246\,
            in2 => \N__44808\,
            in3 => \N__45540\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45368\,
            in1 => \N__45346\,
            in2 => \_gnd_net_\,
            in3 => \N__51315\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51314\,
            in1 => \N__45274\,
            in2 => \_gnd_net_\,
            in3 => \N__45247\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__51313\,
            in1 => \N__41476\,
            in2 => \N__45192\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39579\,
            in1 => \N__44617\,
            in2 => \_gnd_net_\,
            in3 => \N__51316\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39578\,
            in1 => \N__51321\,
            in2 => \_gnd_net_\,
            in3 => \N__44613\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50830\,
            ce => \N__49244\,
            sr => \N__50280\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39560\,
            in1 => \N__51319\,
            in2 => \_gnd_net_\,
            in3 => \N__44807\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50830\,
            ce => \N__49244\,
            sr => \N__50280\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39543\,
            in1 => \N__51320\,
            in2 => \_gnd_net_\,
            in3 => \N__44670\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50830\,
            ce => \N__49244\,
            sr => \N__50280\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39519\,
            in1 => \N__51322\,
            in2 => \_gnd_net_\,
            in3 => \N__48216\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50830\,
            ce => \N__49244\,
            sr => \N__50280\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__41373\,
            in1 => \N__41396\,
            in2 => \N__39489\,
            in3 => \N__39498\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__39497\,
            in1 => \N__41372\,
            in2 => \N__41400\,
            in3 => \N__39485\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48962\,
            in1 => \N__48937\,
            in2 => \_gnd_net_\,
            in3 => \N__51518\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50818\,
            ce => \N__49242\,
            sr => \N__50289\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51517\,
            in1 => \N__47820\,
            in2 => \_gnd_net_\,
            in3 => \N__40932\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50818\,
            ce => \N__49242\,
            sr => \N__50289\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47856\,
            in1 => \N__39472\,
            in2 => \_gnd_net_\,
            in3 => \N__51519\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50818\,
            ce => \N__49242\,
            sr => \N__50289\
        );

    \current_shift_inst.timer_s1.counter_0_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49074\,
            in1 => \N__39445\,
            in2 => \_gnd_net_\,
            in3 => \N__39426\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_1_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49029\,
            in1 => \N__39772\,
            in2 => \_gnd_net_\,
            in3 => \N__39753\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_2_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49075\,
            in1 => \N__39748\,
            in2 => \_gnd_net_\,
            in3 => \N__39732\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_3_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49030\,
            in1 => \N__39727\,
            in2 => \_gnd_net_\,
            in3 => \N__39711\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_4_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49076\,
            in1 => \N__39700\,
            in2 => \_gnd_net_\,
            in3 => \N__39684\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_5_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49031\,
            in1 => \N__39673\,
            in2 => \_gnd_net_\,
            in3 => \N__39657\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_6_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49077\,
            in1 => \N__39652\,
            in2 => \_gnd_net_\,
            in3 => \N__39636\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_7_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49032\,
            in1 => \N__39631\,
            in2 => \_gnd_net_\,
            in3 => \N__39615\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__50809\,
            ce => \N__40314\,
            sr => \N__50297\
        );

    \current_shift_inst.timer_s1.counter_8_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49081\,
            in1 => \N__39604\,
            in2 => \_gnd_net_\,
            in3 => \N__39582\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_9_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49085\,
            in1 => \N__40015\,
            in2 => \_gnd_net_\,
            in3 => \N__39993\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_10_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49078\,
            in1 => \N__39988\,
            in2 => \_gnd_net_\,
            in3 => \N__39972\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_11_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49082\,
            in1 => \N__39967\,
            in2 => \_gnd_net_\,
            in3 => \N__39951\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_12_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49079\,
            in1 => \N__39943\,
            in2 => \_gnd_net_\,
            in3 => \N__39924\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_13_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49083\,
            in1 => \N__39913\,
            in2 => \_gnd_net_\,
            in3 => \N__39897\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_14_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49080\,
            in1 => \N__39886\,
            in2 => \_gnd_net_\,
            in3 => \N__39870\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_15_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49084\,
            in1 => \N__39865\,
            in2 => \_gnd_net_\,
            in3 => \N__39849\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__50801\,
            ce => \N__40322\,
            sr => \N__50304\
        );

    \current_shift_inst.timer_s1.counter_16_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49025\,
            in1 => \N__39841\,
            in2 => \_gnd_net_\,
            in3 => \N__39819\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_17_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49090\,
            in1 => \N__39802\,
            in2 => \_gnd_net_\,
            in3 => \N__40242\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_18_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49026\,
            in1 => \N__40237\,
            in2 => \_gnd_net_\,
            in3 => \N__40221\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_19_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49091\,
            in1 => \N__40216\,
            in2 => \_gnd_net_\,
            in3 => \N__40197\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_20_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49027\,
            in1 => \N__40189\,
            in2 => \_gnd_net_\,
            in3 => \N__40170\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_21_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49092\,
            in1 => \N__40162\,
            in2 => \_gnd_net_\,
            in3 => \N__40143\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_22_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49028\,
            in1 => \N__40132\,
            in2 => \_gnd_net_\,
            in3 => \N__40116\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_23_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49093\,
            in1 => \N__40105\,
            in2 => \_gnd_net_\,
            in3 => \N__40089\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__50793\,
            ce => \N__40315\,
            sr => \N__50313\
        );

    \current_shift_inst.timer_s1.counter_24_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49086\,
            in1 => \N__40081\,
            in2 => \_gnd_net_\,
            in3 => \N__40059\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \current_shift_inst.timer_s1.counter_25_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49094\,
            in1 => \N__40045\,
            in2 => \_gnd_net_\,
            in3 => \N__40029\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \current_shift_inst.timer_s1.counter_26_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49087\,
            in1 => \N__40405\,
            in2 => \_gnd_net_\,
            in3 => \N__40386\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \current_shift_inst.timer_s1.counter_27_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49095\,
            in1 => \N__40381\,
            in2 => \_gnd_net_\,
            in3 => \N__40365\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \current_shift_inst.timer_s1.counter_28_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49088\,
            in1 => \N__40361\,
            in2 => \_gnd_net_\,
            in3 => \N__40347\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \current_shift_inst.timer_s1.counter_29_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__40337\,
            in1 => \N__49089\,
            in2 => \_gnd_net_\,
            in3 => \N__40344\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50783\,
            ce => \N__40323\,
            sr => \N__50320\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__41324\,
            in1 => \N__40280\,
            in2 => \N__40266\,
            in3 => \N__41346\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110001"
        )
    port map (
            in0 => \N__41345\,
            in1 => \N__41323\,
            in2 => \N__40284\,
            in3 => \N__40265\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47894\,
            in1 => \N__40736\,
            in2 => \_gnd_net_\,
            in3 => \N__51501\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51502\,
            in1 => \_gnd_net_\,
            in2 => \N__40251\,
            in3 => \N__47895\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50778\,
            ce => \N__49239\,
            sr => \N__50329\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__42570\,
            in1 => \N__42456\,
            in2 => \_gnd_net_\,
            in3 => \N__46943\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42458\,
            in1 => \N__46936\,
            in2 => \N__46892\,
            in3 => \N__42373\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__42659\,
            in1 => \N__41614\,
            in2 => \N__40428\,
            in3 => \N__42561\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40416\,
            in1 => \N__43855\,
            in2 => \N__40425\,
            in3 => \N__43286\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43512\,
            in1 => \N__42717\,
            in2 => \N__43348\,
            in3 => \N__42776\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011001010"
        )
    port map (
            in0 => \N__46560\,
            in1 => \N__43035\,
            in2 => \N__46764\,
            in3 => \N__46401\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101000"
        )
    port map (
            in0 => \N__42855\,
            in1 => \N__46713\,
            in2 => \N__46421\,
            in3 => \N__46565\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011001010"
        )
    port map (
            in0 => \N__46561\,
            in1 => \N__42924\,
            in2 => \N__46765\,
            in3 => \N__46402\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__46394\,
            in1 => \N__46563\,
            in2 => \N__43488\,
            in3 => \N__46711\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101000"
        )
    port map (
            in0 => \N__42252\,
            in1 => \N__46712\,
            in2 => \N__46420\,
            in3 => \N__46564\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011000101"
        )
    port map (
            in0 => \N__46562\,
            in1 => \N__42327\,
            in2 => \N__46766\,
            in3 => \N__46403\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50769\,
            ce => 'H',
            sr => \N__50351\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__46539\,
            in1 => \N__46778\,
            in2 => \N__43185\,
            in3 => \N__46417\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__46776\,
            in1 => \N__46542\,
            in2 => \N__46424\,
            in3 => \N__43305\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__46538\,
            in1 => \N__46416\,
            in2 => \N__42798\,
            in3 => \N__46779\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__46777\,
            in1 => \N__46543\,
            in2 => \N__46425\,
            in3 => \N__43251\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__46775\,
            in1 => \N__46541\,
            in2 => \N__46423\,
            in3 => \N__43371\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__46774\,
            in1 => \N__46540\,
            in2 => \N__46422\,
            in3 => \N__42741\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50767\,
            ce => 'H',
            sr => \N__50357\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__46388\,
            in1 => \N__46583\,
            in2 => \N__43824\,
            in3 => \N__46762\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__46579\,
            in1 => \N__46390\,
            in2 => \N__46782\,
            in3 => \N__43062\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__46581\,
            in1 => \N__46392\,
            in2 => \N__46784\,
            in3 => \N__43743\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__46389\,
            in1 => \N__46584\,
            in2 => \N__43758\,
            in3 => \N__46763\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__46580\,
            in1 => \N__46391\,
            in2 => \N__46783\,
            in3 => \N__43881\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__46387\,
            in1 => \N__46582\,
            in2 => \N__43131\,
            in3 => \N__46761\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50764\,
            ce => 'H',
            sr => \N__50363\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__46393\,
            in1 => \N__46546\,
            in2 => \N__46785\,
            in3 => \N__43941\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50761\,
            ce => 'H',
            sr => \N__50368\
        );

    \phase_controller_inst1.stoper_hc.time_passed_er_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40517\,
            lcout => \phase_controller_inst1.stoper_hc.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50909\,
            ce => \N__40437\,
            sr => \N__50231\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__48711\,
            in1 => \N__40587\,
            in2 => \_gnd_net_\,
            in3 => \N__40574\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50903\,
            ce => 'H',
            sr => \N__50234\
        );

    \phase_controller_inst1.stoper_hc.running_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__40516\,
            in1 => \N__40486\,
            in2 => \_gnd_net_\,
            in3 => \N__40446\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50903\,
            ce => 'H',
            sr => \N__50234\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_30_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101011101"
        )
    port map (
            in0 => \N__40553\,
            in1 => \N__40518\,
            in2 => \N__40488\,
            in3 => \N__40464\,
            lcout => \phase_controller_inst1.stoper_hc.N_46\,
            ltout => \phase_controller_inst1.stoper_hc.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_sbtinv_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40440\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.N_46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__40760\,
            in1 => \N__44169\,
            in2 => \N__40796\,
            in3 => \N__40818\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__40817\,
            in1 => \N__40761\,
            in2 => \N__40797\,
            in3 => \N__44168\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45471\,
            in1 => \N__51440\,
            in2 => \_gnd_net_\,
            in3 => \N__45501\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50891\,
            ce => \N__48852\,
            sr => \N__50241\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47999\,
            in1 => \N__51441\,
            in2 => \_gnd_net_\,
            in3 => \N__48037\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50891\,
            ce => \N__48852\,
            sr => \N__50241\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51437\,
            in1 => \N__47888\,
            in2 => \_gnd_net_\,
            in3 => \N__40746\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50891\,
            ce => \N__48852\,
            sr => \N__50241\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48308\,
            in1 => \N__51439\,
            in2 => \_gnd_net_\,
            in3 => \N__48284\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50891\,
            ce => \N__48852\,
            sr => \N__50241\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51438\,
            in1 => \N__47818\,
            in2 => \_gnd_net_\,
            in3 => \N__40924\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50891\,
            ce => \N__48852\,
            sr => \N__50241\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__44037\,
            in1 => \N__40941\,
            in2 => \N__40692\,
            in3 => \N__40669\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__40940\,
            in1 => \N__40690\,
            in2 => \N__40671\,
            in3 => \N__44036\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51436\,
            in1 => \N__41483\,
            in2 => \_gnd_net_\,
            in3 => \N__45190\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50884\,
            ce => \N__48812\,
            sr => \N__50246\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40928\,
            in1 => \N__47817\,
            in2 => \_gnd_net_\,
            in3 => \N__51435\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__40896\,
            in1 => \N__40887\,
            in2 => \N__47955\,
            in3 => \N__40866\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__51762\,
            in1 => \N__51723\,
            in2 => \N__51460\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50874\,
            ce => \N__48853\,
            sr => \N__50250\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__40895\,
            in1 => \N__40886\,
            in2 => \N__47954\,
            in3 => \N__40865\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41160\,
            in1 => \N__44929\,
            in2 => \_gnd_net_\,
            in3 => \N__40836\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41177\,
            in1 => \N__48109\,
            in2 => \_gnd_net_\,
            in3 => \N__40833\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41161\,
            in1 => \N__44324\,
            in2 => \_gnd_net_\,
            in3 => \N__40830\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41178\,
            in1 => \N__44300\,
            in2 => \_gnd_net_\,
            in3 => \N__40827\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41162\,
            in1 => \N__44276\,
            in2 => \_gnd_net_\,
            in3 => \N__40968\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41179\,
            in1 => \N__44252\,
            in2 => \_gnd_net_\,
            in3 => \N__40965\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41163\,
            in1 => \N__44228\,
            in2 => \_gnd_net_\,
            in3 => \N__40962\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41180\,
            in1 => \N__44570\,
            in2 => \_gnd_net_\,
            in3 => \N__40959\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__50865\,
            ce => \N__41049\,
            sr => \N__50258\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41159\,
            in1 => \N__44546\,
            in2 => \_gnd_net_\,
            in3 => \N__40956\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41167\,
            in1 => \N__44522\,
            in2 => \_gnd_net_\,
            in3 => \N__40953\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41156\,
            in1 => \N__44498\,
            in2 => \_gnd_net_\,
            in3 => \N__40950\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41164\,
            in1 => \N__44441\,
            in2 => \_gnd_net_\,
            in3 => \N__40947\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41157\,
            in1 => \N__44417\,
            in2 => \_gnd_net_\,
            in3 => \N__40944\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41165\,
            in1 => \N__44393\,
            in2 => \_gnd_net_\,
            in3 => \N__40995\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41158\,
            in1 => \N__44369\,
            in2 => \_gnd_net_\,
            in3 => \N__40992\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41166\,
            in1 => \N__44873\,
            in2 => \_gnd_net_\,
            in3 => \N__40989\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__50852\,
            ce => \N__41048\,
            sr => \N__50266\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41152\,
            in1 => \N__44849\,
            in2 => \_gnd_net_\,
            in3 => \N__40986\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41181\,
            in1 => \N__44825\,
            in2 => \_gnd_net_\,
            in3 => \N__40983\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41153\,
            in1 => \N__44768\,
            in2 => \_gnd_net_\,
            in3 => \N__40980\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41182\,
            in1 => \N__44744\,
            in2 => \_gnd_net_\,
            in3 => \N__40977\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41154\,
            in1 => \N__44720\,
            in2 => \_gnd_net_\,
            in3 => \N__40974\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41183\,
            in1 => \N__44696\,
            in2 => \_gnd_net_\,
            in3 => \N__40971\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41155\,
            in1 => \N__44636\,
            in2 => \_gnd_net_\,
            in3 => \N__41205\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41184\,
            in1 => \N__45209\,
            in2 => \_gnd_net_\,
            in3 => \N__41202\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__50842\,
            ce => \N__41041\,
            sr => \N__50272\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41137\,
            in1 => \N__45134\,
            in2 => \_gnd_net_\,
            in3 => \N__41199\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41141\,
            in1 => \N__45110\,
            in2 => \_gnd_net_\,
            in3 => \N__41196\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41138\,
            in1 => \N__45074\,
            in2 => \_gnd_net_\,
            in3 => \N__41193\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41142\,
            in1 => \N__45002\,
            in2 => \_gnd_net_\,
            in3 => \N__41190\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41139\,
            in1 => \N__45090\,
            in2 => \_gnd_net_\,
            in3 => \N__41187\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__45018\,
            in1 => \N__41140\,
            in2 => \_gnd_net_\,
            in3 => \N__41052\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50831\,
            ce => \N__41040\,
            sr => \N__50281\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46980\,
            in2 => \N__41243\,
            in3 => \N__46995\,
            lcout => \phase_controller_inst2.stoper_hc.N_265_i\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47155\,
            in1 => \N__45749\,
            in2 => \_gnd_net_\,
            in3 => \N__41247\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__47144\,
            in1 => \N__45722\,
            in2 => \N__41244\,
            in3 => \N__41229\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47156\,
            in1 => \N__45692\,
            in2 => \_gnd_net_\,
            in3 => \N__41226\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47145\,
            in1 => \N__45668\,
            in2 => \_gnd_net_\,
            in3 => \N__41223\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47157\,
            in1 => \N__45617\,
            in2 => \_gnd_net_\,
            in3 => \N__41220\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47146\,
            in1 => \N__45581\,
            in2 => \_gnd_net_\,
            in3 => \N__41217\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47158\,
            in1 => \N__45995\,
            in2 => \_gnd_net_\,
            in3 => \N__41214\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50819\,
            ce => 'H',
            sr => \N__50290\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47165\,
            in1 => \N__45968\,
            in2 => \_gnd_net_\,
            in3 => \N__41211\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47140\,
            in1 => \N__45947\,
            in2 => \_gnd_net_\,
            in3 => \N__41208\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47162\,
            in1 => \N__45923\,
            in2 => \_gnd_net_\,
            in3 => \N__41274\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47141\,
            in1 => \N__45887\,
            in2 => \_gnd_net_\,
            in3 => \N__41271\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__45860\,
            in2 => \_gnd_net_\,
            in3 => \N__41268\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47142\,
            in1 => \N__45824\,
            in2 => \_gnd_net_\,
            in3 => \N__41265\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47164\,
            in1 => \N__45779\,
            in2 => \_gnd_net_\,
            in3 => \N__41262\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47143\,
            in1 => \N__44913\,
            in2 => \_gnd_net_\,
            in3 => \N__41259\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__50810\,
            ce => 'H',
            sr => \N__50298\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47147\,
            in1 => \N__44893\,
            in2 => \_gnd_net_\,
            in3 => \N__41256\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47133\,
            in1 => \N__45294\,
            in2 => \_gnd_net_\,
            in3 => \N__41253\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47148\,
            in1 => \N__45311\,
            in2 => \_gnd_net_\,
            in3 => \N__41250\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47134\,
            in1 => \N__41390\,
            in2 => \_gnd_net_\,
            in3 => \N__41376\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47149\,
            in1 => \N__41371\,
            in2 => \_gnd_net_\,
            in3 => \N__41355\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47135\,
            in1 => \N__51013\,
            in2 => \_gnd_net_\,
            in3 => \N__41352\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47150\,
            in1 => \N__51043\,
            in2 => \_gnd_net_\,
            in3 => \N__41349\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47136\,
            in1 => \N__41344\,
            in2 => \_gnd_net_\,
            in3 => \N__41328\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__50802\,
            ce => 'H',
            sr => \N__50305\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47151\,
            in1 => \N__41325\,
            in2 => \_gnd_net_\,
            in3 => \N__41310\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47159\,
            in1 => \N__41499\,
            in2 => \_gnd_net_\,
            in3 => \N__41307\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47152\,
            in1 => \N__41516\,
            in2 => \_gnd_net_\,
            in3 => \N__41304\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47160\,
            in1 => \N__41291\,
            in2 => \_gnd_net_\,
            in3 => \N__41277\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47153\,
            in1 => \N__41540\,
            in2 => \_gnd_net_\,
            in3 => \N__41526\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47161\,
            in1 => \N__41415\,
            in2 => \_gnd_net_\,
            in3 => \N__41523\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47154\,
            in1 => \N__41444\,
            in2 => \_gnd_net_\,
            in3 => \N__41520\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50794\,
            ce => 'H',
            sr => \N__50314\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__41498\,
            in1 => \N__49337\,
            in2 => \N__41517\,
            in3 => \N__41454\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__41453\,
            in1 => \N__41515\,
            in2 => \N__49341\,
            in3 => \N__41497\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41484\,
            in1 => \N__45191\,
            in2 => \_gnd_net_\,
            in3 => \N__51622\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50784\,
            ce => \N__49240\,
            sr => \N__50321\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49205\,
            in1 => \N__49154\,
            in2 => \_gnd_net_\,
            in3 => \N__51623\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50784\,
            ce => \N__49240\,
            sr => \N__50321\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011111101"
        )
    port map (
            in0 => \N__41413\,
            in1 => \N__42170\,
            in2 => \N__41445\,
            in3 => \N__41423\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__42171\,
            in1 => \N__41440\,
            in2 => \N__41427\,
            in3 => \N__41414\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51621\,
            in1 => \N__42198\,
            in2 => \_gnd_net_\,
            in3 => \N__44984\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50784\,
            ce => \N__49240\,
            sr => \N__50321\
        );

    \phase_controller_inst2.start_timer_hc_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__41925\,
            in1 => \N__42005\,
            in2 => \N__42162\,
            in3 => \N__42128\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50779\,
            ce => \N__43641\,
            sr => \N__50330\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0_30_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__42003\,
            in1 => \N__42089\,
            in2 => \N__42068\,
            in3 => \N__47174\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_30_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011111111"
        )
    port map (
            in0 => \N__42090\,
            in1 => \N__42064\,
            in2 => \N__47178\,
            in3 => \N__42004\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__41819\,
            in1 => \N__41961\,
            in2 => \N__41946\,
            in3 => \N__41924\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50779\,
            ce => \N__43641\,
            sr => \N__50330\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41790\,
            in2 => \N__41738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41693\,
            in2 => \N__41664\,
            in3 => \N__41634\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41613\,
            in2 => \N__41586\,
            in3 => \N__41556\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42655\,
            in2 => \N__42618\,
            in3 => \N__42585\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42582\,
            in2 => \N__42569\,
            in3 => \N__42507\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46872\,
            in2 => \N__42504\,
            in3 => \N__42486\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46932\,
            in2 => \N__42483\,
            in3 => \N__42465\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42457\,
            in2 => \N__42420\,
            in3 => \N__42387\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42369\,
            in2 => \N__42345\,
            in3 => \N__42321\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42292\,
            in2 => \N__42273\,
            in3 => \N__42246\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42222\,
            in2 => \N__43053\,
            in3 => \N__43029\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46806\,
            in2 => \N__43026\,
            in3 => \N__43008\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46219\,
            in2 => \N__43005\,
            in3 => \N__42987\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42959\,
            in2 => \N__42942\,
            in3 => \N__42918\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42892\,
            in2 => \N__42873\,
            in3 => \N__42849\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42825\,
            in2 => \N__46167\,
            in3 => \N__42789\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42762\,
            in2 => \N__47451\,
            in3 => \N__42735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42718\,
            in2 => \N__47406\,
            in3 => \N__42672\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43513\,
            in2 => \N__47358\,
            in3 => \N__43476\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43461\,
            in2 => \N__47328\,
            in3 => \N__43416\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43395\,
            in2 => \N__47298\,
            in3 => \N__43365\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43335\,
            in2 => \N__47271\,
            in3 => \N__43299\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43272\,
            in2 => \N__47241\,
            in3 => \N__43245\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43218\,
            in2 => \N__47211\,
            in3 => \N__43176\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43155\,
            in2 => \N__47748\,
            in3 => \N__43119\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43092\,
            in2 => \N__47712\,
            in3 => \N__43056\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47682\,
            in2 => \N__43977\,
            in3 => \N__43935\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43905\,
            in2 => \N__47652\,
            in3 => \N__43875\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43842\,
            in2 => \N__47625\,
            in3 => \N__43815\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43785\,
            in2 => \N__47514\,
            in3 => \N__43749\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46516\,
            in1 => \N__47499\,
            in2 => \N__43716\,
            in3 => \N__43746\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47607\,
            in2 => \_gnd_net_\,
            in3 => \N__43737\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_5_LC_17_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \phase_controller_inst1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50752\,
            ce => \N__43669\,
            sr => \N__50384\
        );

    \phase_controller_inst1.test_LC_17_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43700\,
            in2 => \_gnd_net_\,
            in3 => \N__43707\,
            lcout => test_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50752\,
            ce => \N__43669\,
            sr => \N__50384\
        );

    \phase_controller_inst2.stoper_tr.time_passed_er_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44127\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50910\,
            ce => \N__44046\,
            sr => \N__50232\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45543\,
            in1 => \N__45561\,
            in2 => \_gnd_net_\,
            in3 => \N__51446\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50904\,
            ce => \N__48867\,
            sr => \N__50235\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51445\,
            in1 => \N__48459\,
            in2 => \_gnd_net_\,
            in3 => \N__48429\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50904\,
            ce => \N__48867\,
            sr => \N__50235\
        );

    \phase_controller_inst2.stoper_tr.running_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__44145\,
            in1 => \N__44074\,
            in2 => \_gnd_net_\,
            in3 => \N__44058\,
            lcout => \phase_controller_inst2.running\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50898\,
            ce => 'H',
            sr => \N__50238\
        );

    \phase_controller_inst2.stoper_tr.time_passed_sbtinv_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44057\,
            lcout => \phase_controller_inst2.stoper_tr.N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51442\,
            in1 => \N__51693\,
            in2 => \_gnd_net_\,
            in3 => \N__51654\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50892\,
            ce => \N__48824\,
            sr => \N__50242\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51443\,
            in1 => \N__48597\,
            in2 => \_gnd_net_\,
            in3 => \N__48567\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50892\,
            ce => \N__48824\,
            sr => \N__50242\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49380\,
            in1 => \N__49421\,
            in2 => \_gnd_net_\,
            in3 => \N__51444\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50892\,
            ce => \N__48824\,
            sr => \N__50242\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45345\,
            in1 => \N__45415\,
            in2 => \N__44479\,
            in3 => \N__45462\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__51431\,
            in1 => \N__44345\,
            in2 => \N__44480\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44475\,
            in2 => \N__44334\,
            in3 => \N__51432\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50885\,
            ce => \N__49251\,
            sr => \N__50247\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44323\,
            in2 => \N__44936\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44299\,
            in2 => \N__48116\,
            in3 => \N__44331\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44275\,
            in2 => \N__44328\,
            in3 => \N__44307\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44251\,
            in2 => \N__44304\,
            in3 => \N__44283\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44227\,
            in2 => \N__44280\,
            in3 => \N__44259\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44569\,
            in2 => \N__44256\,
            in3 => \N__44235\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44545\,
            in2 => \N__44232\,
            in3 => \N__44211\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44521\,
            in2 => \N__44574\,
            in3 => \N__44553\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__50875\,
            ce => \N__48089\,
            sr => \N__50251\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44497\,
            in2 => \N__44550\,
            in3 => \N__44529\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44440\,
            in2 => \N__44526\,
            in3 => \N__44505\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44416\,
            in2 => \N__44502\,
            in3 => \N__44448\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44392\,
            in2 => \N__44445\,
            in3 => \N__44424\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44368\,
            in2 => \N__44421\,
            in3 => \N__44400\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44872\,
            in2 => \N__44397\,
            in3 => \N__44376\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44848\,
            in2 => \N__44373\,
            in3 => \N__44352\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44824\,
            in2 => \N__44877\,
            in3 => \N__44856\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__50866\,
            ce => \N__48088\,
            sr => \N__50259\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44767\,
            in2 => \N__44853\,
            in3 => \N__44832\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44743\,
            in2 => \N__44829\,
            in3 => \N__44775\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44719\,
            in2 => \N__44772\,
            in3 => \N__44751\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44695\,
            in2 => \N__44748\,
            in3 => \N__44727\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44635\,
            in2 => \N__44724\,
            in3 => \N__44703\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45208\,
            in2 => \N__44700\,
            in3 => \N__44643\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45133\,
            in2 => \N__44640\,
            in3 => \N__44577\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45109\,
            in2 => \N__45213\,
            in3 => \N__45141\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__50853\,
            ce => \N__48087\,
            sr => \N__50267\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45073\,
            in2 => \N__45138\,
            in3 => \N__45117\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45001\,
            in2 => \N__45114\,
            in3 => \N__45093\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45089\,
            in2 => \N__45078\,
            in3 => \N__45021\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45017\,
            in2 => \N__45006\,
            in3 => \N__44946\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44943\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44940\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50843\,
            ce => \N__48074\,
            sr => \N__50273\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__44911\,
            in1 => \N__44894\,
            in2 => \N__45513\,
            in3 => \N__45435\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__45434\,
            in1 => \N__44912\,
            in2 => \N__44898\,
            in3 => \N__45509\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45541\,
            in1 => \N__45557\,
            in2 => \_gnd_net_\,
            in3 => \N__51600\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51603\,
            in1 => \_gnd_net_\,
            in2 => \N__45546\,
            in3 => \N__45542\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50832\,
            ce => \N__49245\,
            sr => \N__50282\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51602\,
            in1 => \N__45500\,
            in2 => \_gnd_net_\,
            in3 => \N__45466\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50832\,
            ce => \N__49245\,
            sr => \N__50282\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45424\,
            in1 => \N__45393\,
            in2 => \_gnd_net_\,
            in3 => \N__51604\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50832\,
            ce => \N__49245\,
            sr => \N__50282\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51601\,
            in1 => \N__45372\,
            in2 => \_gnd_net_\,
            in3 => \N__45348\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50832\,
            ce => \N__49245\,
            sr => \N__50282\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__45293\,
            in1 => \N__45222\,
            in2 => \N__49440\,
            in3 => \N__45310\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__49439\,
            in2 => \N__45312\,
            in3 => \N__45292\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__45279\,
            in1 => \N__45251\,
            in2 => \N__51624\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50820\,
            ce => \N__49243\,
            sr => \N__50291\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48036\,
            in1 => \N__51612\,
            in2 => \_gnd_net_\,
            in3 => \N__48003\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50820\,
            ce => \N__49243\,
            sr => \N__50291\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49350\,
            in2 => \N__45765\,
            in3 => \N__46976\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48471\,
            in2 => \N__45735\,
            in3 => \N__45753\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45708\,
            in2 => \N__48399\,
            in3 => \N__45726\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45702\,
            in2 => \N__45678\,
            in3 => \N__45696\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45669\,
            in1 => \N__45654\,
            in2 => \N__45642\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45603\,
            in2 => \N__45633\,
            in3 => \N__45618\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45567\,
            in2 => \N__45597\,
            in3 => \N__45582\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45996\,
            in1 => \N__48537\,
            in2 => \N__45981\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45954\,
            in2 => \N__48327\,
            in3 => \N__45972\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45933\,
            in2 => \N__48246\,
            in3 => \N__45948\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49263\,
            in2 => \N__45909\,
            in3 => \N__45927\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45900\,
            in2 => \N__45873\,
            in3 => \N__45888\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45861\,
            in1 => \N__45831\,
            in2 => \N__45846\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45825\,
            in1 => \N__45810\,
            in2 => \N__45801\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45789\,
            in2 => \N__46158\,
            in3 => \N__45780\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46149\,
            in2 => \N__46137\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46122\,
            in2 => \N__46113\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46098\,
            in2 => \N__46083\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48231\,
            in2 => \N__50985\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46065\,
            in2 => \N__46056\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46044\,
            in2 => \N__46038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46029\,
            in2 => \N__46017\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47199\,
            in2 => \N__47193\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_0_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_LUT4_0_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47181\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__47107\,
            in1 => \N__46994\,
            in2 => \_gnd_net_\,
            in3 => \N__46975\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50785\,
            ce => 'H',
            sr => \N__50322\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__46719\,
            in1 => \N__46596\,
            in2 => \N__46419\,
            in3 => \N__46956\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50780\,
            ce => 'H',
            sr => \N__50331\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__46595\,
            in1 => \N__46383\,
            in2 => \N__46908\,
            in3 => \N__46720\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50780\,
            ce => 'H',
            sr => \N__50331\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__46593\,
            in1 => \N__46384\,
            in2 => \N__46848\,
            in3 => \N__46768\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50773\,
            ce => 'H',
            sr => \N__50337\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__46767\,
            in1 => \N__46594\,
            in2 => \N__46434\,
            in3 => \N__46385\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50773\,
            ce => 'H',
            sr => \N__50337\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46203\,
            in2 => \N__46185\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47487\,
            in2 => \N__47469\,
            in3 => \N__47442\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47439\,
            in2 => \N__47424\,
            in3 => \N__47397\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47394\,
            in2 => \N__47376\,
            in3 => \N__47349\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47346\,
            in2 => \N__47608\,
            in3 => \N__47316\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47313\,
            in2 => \N__47610\,
            in3 => \N__47289\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47286\,
            in2 => \N__47609\,
            in3 => \N__47262\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47590\,
            in2 => \N__47259\,
            in3 => \N__47232\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47594\,
            in2 => \N__47229\,
            in3 => \N__47202\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47766\,
            in2 => \N__47611\,
            in3 => \N__47736\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47598\,
            in2 => \N__47733\,
            in3 => \N__47703\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47700\,
            in2 => \N__47612\,
            in3 => \N__47676\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47602\,
            in2 => \N__47673\,
            in3 => \N__47643\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47640\,
            in2 => \N__47613\,
            in3 => \N__47616\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47606\,
            in2 => \N__47535\,
            in3 => \N__47505\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47502\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48501\,
            in1 => \N__48525\,
            in2 => \_gnd_net_\,
            in3 => \N__51620\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50912\,
            ce => \N__48861\,
            sr => \N__50236\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51616\,
            in1 => \N__48307\,
            in2 => \_gnd_net_\,
            in3 => \N__48283\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48382\,
            in1 => \N__48338\,
            in2 => \_gnd_net_\,
            in3 => \N__51617\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51618\,
            in1 => \_gnd_net_\,
            in2 => \N__47922\,
            in3 => \N__48383\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50911\,
            ce => \N__48875\,
            sr => \N__50239\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49318\,
            in1 => \N__49301\,
            in2 => \_gnd_net_\,
            in3 => \N__51619\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50906\,
            ce => \N__48860\,
            sr => \N__50243\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48454\,
            in1 => \N__48431\,
            in2 => \_gnd_net_\,
            in3 => \N__51430\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49296\,
            in1 => \N__48282\,
            in2 => \N__48384\,
            in3 => \N__47887\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__47854\,
            in1 => \N__47819\,
            in2 => \N__47784\,
            in3 => \N__48177\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49297\,
            in1 => \N__51433\,
            in2 => \_gnd_net_\,
            in3 => \N__49322\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48571\,
            in2 => \_gnd_net_\,
            in3 => \N__48213\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48430\,
            in1 => \N__48492\,
            in2 => \N__49425\,
            in3 => \N__48038\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48162\,
            in2 => \N__48129\,
            in3 => \N__51694\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48572\,
            in1 => \N__51434\,
            in2 => \_gnd_net_\,
            in3 => \N__48592\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48117\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50893\,
            ce => \N__48093\,
            sr => \N__50252\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48523\,
            in1 => \N__48493\,
            in2 => \_gnd_net_\,
            in3 => \N__51581\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47992\,
            in1 => \N__48039\,
            in2 => \_gnd_net_\,
            in3 => \N__51580\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49476\,
            in1 => \N__49497\,
            in2 => \_gnd_net_\,
            in3 => \N__51595\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50886\,
            ce => \N__48868\,
            sr => \N__50260\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51087\,
            in1 => \N__51127\,
            in2 => \_gnd_net_\,
            in3 => \N__51596\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50886\,
            ce => \N__48868\,
            sr => \N__50260\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51593\,
            in1 => \N__48593\,
            in2 => \_gnd_net_\,
            in3 => \N__48573\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50876\,
            ce => \N__49250\,
            sr => \N__50268\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48524\,
            in1 => \N__51594\,
            in2 => \_gnd_net_\,
            in3 => \N__48500\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50876\,
            ce => \N__49250\,
            sr => \N__50268\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51592\,
            in1 => \N__48455\,
            in2 => \_gnd_net_\,
            in3 => \N__48432\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50876\,
            ce => \N__49250\,
            sr => \N__50268\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51556\,
            in1 => \N__51082\,
            in2 => \_gnd_net_\,
            in3 => \N__51128\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50867\,
            ce => \N__49249\,
            sr => \N__50274\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__51716\,
            in1 => \N__51555\,
            in2 => \_gnd_net_\,
            in3 => \N__51765\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50867\,
            ce => \N__49249\,
            sr => \N__50274\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51557\,
            in1 => \N__48381\,
            in2 => \_gnd_net_\,
            in3 => \N__48345\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50867\,
            ce => \N__49249\,
            sr => \N__50274\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48312\,
            in1 => \N__48285\,
            in2 => \_gnd_net_\,
            in3 => \N__51558\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50867\,
            ce => \N__49249\,
            sr => \N__50274\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__51065\,
            in1 => \N__51050\,
            in2 => \N__51027\,
            in3 => \N__50996\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__49496\,
            in1 => \N__49474\,
            in2 => \N__51579\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49419\,
            in1 => \N__51522\,
            in2 => \_gnd_net_\,
            in3 => \N__49372\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49492\,
            in1 => \N__49475\,
            in2 => \_gnd_net_\,
            in3 => \N__51554\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50844\,
            ce => \N__49247\,
            sr => \N__50292\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49420\,
            in1 => \N__51551\,
            in2 => \_gnd_net_\,
            in3 => \N__49373\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50833\,
            ce => \N__49246\,
            sr => \N__50299\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51552\,
            in1 => \N__51696\,
            in2 => \_gnd_net_\,
            in3 => \N__51653\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50833\,
            ce => \N__49246\,
            sr => \N__50299\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49323\,
            in1 => \N__49302\,
            in2 => \_gnd_net_\,
            in3 => \N__51553\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50833\,
            ce => \N__49246\,
            sr => \N__50299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49153\,
            in1 => \N__49206\,
            in2 => \_gnd_net_\,
            in3 => \N__51521\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49131\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51515\,
            in1 => \N__48963\,
            in2 => \_gnd_net_\,
            in3 => \N__48938\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50899\,
            ce => \N__48876\,
            sr => \N__50261\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51715\,
            in1 => \N__51764\,
            in2 => \_gnd_net_\,
            in3 => \N__51503\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51504\,
            in1 => \N__51695\,
            in2 => \_gnd_net_\,
            in3 => \N__51646\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51559\,
            in1 => \N__51086\,
            in2 => \_gnd_net_\,
            in3 => \N__51129\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__51066\,
            in1 => \N__51054\,
            in2 => \N__51026\,
            in3 => \N__50997\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50966\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50834\,
            ce => 'H',
            sr => \N__50315\
        );

    \CONSTANT_ONE_LUT4_LC_22_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
