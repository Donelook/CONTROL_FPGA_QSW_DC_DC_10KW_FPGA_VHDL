// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Nov 29 2024 16:50:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    test,
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    test22,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output test;
    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output test22;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50662;
    wire N__50661;
    wire N__50660;
    wire N__50651;
    wire N__50650;
    wire N__50649;
    wire N__50642;
    wire N__50641;
    wire N__50640;
    wire N__50633;
    wire N__50632;
    wire N__50631;
    wire N__50624;
    wire N__50623;
    wire N__50622;
    wire N__50615;
    wire N__50614;
    wire N__50613;
    wire N__50606;
    wire N__50605;
    wire N__50604;
    wire N__50597;
    wire N__50596;
    wire N__50595;
    wire N__50588;
    wire N__50587;
    wire N__50586;
    wire N__50579;
    wire N__50578;
    wire N__50577;
    wire N__50570;
    wire N__50569;
    wire N__50568;
    wire N__50561;
    wire N__50560;
    wire N__50559;
    wire N__50552;
    wire N__50551;
    wire N__50550;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50534;
    wire N__50533;
    wire N__50532;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50506;
    wire N__50505;
    wire N__50502;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50489;
    wire N__50484;
    wire N__50481;
    wire N__50476;
    wire N__50473;
    wire N__50472;
    wire N__50469;
    wire N__50468;
    wire N__50465;
    wire N__50460;
    wire N__50457;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50442;
    wire N__50441;
    wire N__50434;
    wire N__50431;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50416;
    wire N__50413;
    wire N__50412;
    wire N__50409;
    wire N__50406;
    wire N__50405;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50380;
    wire N__50377;
    wire N__50376;
    wire N__50375;
    wire N__50372;
    wire N__50367;
    wire N__50364;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50352;
    wire N__50349;
    wire N__50346;
    wire N__50345;
    wire N__50340;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50326;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50318;
    wire N__50313;
    wire N__50310;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50294;
    wire N__50291;
    wire N__50288;
    wire N__50283;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50269;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50261;
    wire N__50258;
    wire N__50255;
    wire N__50252;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50239;
    wire N__50238;
    wire N__50237;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50225;
    wire N__50222;
    wire N__50219;
    wire N__50210;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50192;
    wire N__50189;
    wire N__50184;
    wire N__50179;
    wire N__50178;
    wire N__50175;
    wire N__50174;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50162;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50146;
    wire N__50143;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50125;
    wire N__50124;
    wire N__50123;
    wire N__50122;
    wire N__50121;
    wire N__50118;
    wire N__50115;
    wire N__50110;
    wire N__50107;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50091;
    wire N__50088;
    wire N__50083;
    wire N__50082;
    wire N__50081;
    wire N__50080;
    wire N__50079;
    wire N__50078;
    wire N__50069;
    wire N__50064;
    wire N__50063;
    wire N__50058;
    wire N__50055;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50040;
    wire N__50039;
    wire N__50036;
    wire N__50031;
    wire N__50028;
    wire N__50023;
    wire N__50020;
    wire N__50019;
    wire N__50018;
    wire N__50017;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50013;
    wire N__50012;
    wire N__50011;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50004;
    wire N__50003;
    wire N__50002;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49998;
    wire N__49997;
    wire N__49996;
    wire N__49995;
    wire N__49994;
    wire N__49993;
    wire N__49992;
    wire N__49991;
    wire N__49990;
    wire N__49989;
    wire N__49988;
    wire N__49987;
    wire N__49986;
    wire N__49985;
    wire N__49984;
    wire N__49983;
    wire N__49982;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49976;
    wire N__49975;
    wire N__49974;
    wire N__49973;
    wire N__49972;
    wire N__49971;
    wire N__49970;
    wire N__49969;
    wire N__49968;
    wire N__49967;
    wire N__49966;
    wire N__49965;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49961;
    wire N__49960;
    wire N__49959;
    wire N__49958;
    wire N__49957;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49933;
    wire N__49932;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49926;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49914;
    wire N__49913;
    wire N__49912;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49907;
    wire N__49906;
    wire N__49905;
    wire N__49904;
    wire N__49903;
    wire N__49902;
    wire N__49901;
    wire N__49900;
    wire N__49899;
    wire N__49898;
    wire N__49897;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49558;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49543;
    wire N__49540;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49530;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49519;
    wire N__49518;
    wire N__49517;
    wire N__49516;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49512;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49492;
    wire N__49491;
    wire N__49490;
    wire N__49489;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49478;
    wire N__49477;
    wire N__49476;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49466;
    wire N__49465;
    wire N__49464;
    wire N__49463;
    wire N__49462;
    wire N__49461;
    wire N__49460;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49401;
    wire N__49400;
    wire N__49399;
    wire N__49398;
    wire N__49397;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49393;
    wire N__49392;
    wire N__49391;
    wire N__49390;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49386;
    wire N__49385;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49374;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49047;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49043;
    wire N__49042;
    wire N__49041;
    wire N__49038;
    wire N__49023;
    wire N__49018;
    wire N__49017;
    wire N__49016;
    wire N__49013;
    wire N__49008;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48954;
    wire N__48951;
    wire N__48948;
    wire N__48945;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48928;
    wire N__48925;
    wire N__48924;
    wire N__48923;
    wire N__48920;
    wire N__48917;
    wire N__48914;
    wire N__48911;
    wire N__48908;
    wire N__48905;
    wire N__48898;
    wire N__48897;
    wire N__48894;
    wire N__48891;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48872;
    wire N__48869;
    wire N__48866;
    wire N__48863;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48851;
    wire N__48848;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48832;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48819;
    wire N__48816;
    wire N__48813;
    wire N__48810;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48787;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48775;
    wire N__48774;
    wire N__48773;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48761;
    wire N__48758;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48743;
    wire N__48740;
    wire N__48737;
    wire N__48734;
    wire N__48731;
    wire N__48728;
    wire N__48721;
    wire N__48720;
    wire N__48717;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48698;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48684;
    wire N__48683;
    wire N__48680;
    wire N__48675;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48648;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48613;
    wire N__48608;
    wire N__48605;
    wire N__48602;
    wire N__48599;
    wire N__48596;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48580;
    wire N__48579;
    wire N__48574;
    wire N__48571;
    wire N__48570;
    wire N__48567;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48522;
    wire N__48517;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48494;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48482;
    wire N__48479;
    wire N__48476;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48455;
    wire N__48452;
    wire N__48449;
    wire N__48446;
    wire N__48443;
    wire N__48436;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48428;
    wire N__48425;
    wire N__48422;
    wire N__48421;
    wire N__48414;
    wire N__48411;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48390;
    wire N__48389;
    wire N__48386;
    wire N__48385;
    wire N__48384;
    wire N__48383;
    wire N__48382;
    wire N__48375;
    wire N__48366;
    wire N__48363;
    wire N__48362;
    wire N__48359;
    wire N__48358;
    wire N__48357;
    wire N__48356;
    wire N__48355;
    wire N__48354;
    wire N__48353;
    wire N__48352;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48339;
    wire N__48332;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48328;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48321;
    wire N__48320;
    wire N__48319;
    wire N__48318;
    wire N__48317;
    wire N__48316;
    wire N__48315;
    wire N__48310;
    wire N__48303;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48297;
    wire N__48288;
    wire N__48285;
    wire N__48284;
    wire N__48283;
    wire N__48282;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48275;
    wire N__48274;
    wire N__48273;
    wire N__48272;
    wire N__48271;
    wire N__48270;
    wire N__48269;
    wire N__48268;
    wire N__48267;
    wire N__48260;
    wire N__48257;
    wire N__48252;
    wire N__48247;
    wire N__48244;
    wire N__48243;
    wire N__48242;
    wire N__48239;
    wire N__48224;
    wire N__48223;
    wire N__48222;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48183;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48169;
    wire N__48168;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48163;
    wire N__48162;
    wire N__48161;
    wire N__48160;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48149;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48126;
    wire N__48119;
    wire N__48114;
    wire N__48111;
    wire N__48106;
    wire N__48101;
    wire N__48096;
    wire N__48089;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48061;
    wire N__48056;
    wire N__48049;
    wire N__48044;
    wire N__48035;
    wire N__48032;
    wire N__48017;
    wire N__48014;
    wire N__48007;
    wire N__48004;
    wire N__47999;
    wire N__47996;
    wire N__47985;
    wire N__47980;
    wire N__47961;
    wire N__47932;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47920;
    wire N__47919;
    wire N__47918;
    wire N__47917;
    wire N__47916;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47911;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47871;
    wire N__47868;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47835;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47813;
    wire N__47808;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47775;
    wire N__47770;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47755;
    wire N__47754;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47742;
    wire N__47737;
    wire N__47734;
    wire N__47731;
    wire N__47728;
    wire N__47725;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47695;
    wire N__47694;
    wire N__47693;
    wire N__47690;
    wire N__47689;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47651;
    wire N__47648;
    wire N__47641;
    wire N__47640;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47625;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47602;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47594;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47561;
    wire N__47554;
    wire N__47553;
    wire N__47548;
    wire N__47545;
    wire N__47544;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47524;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47510;
    wire N__47507;
    wire N__47500;
    wire N__47497;
    wire N__47496;
    wire N__47493;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47460;
    wire N__47455;
    wire N__47452;
    wire N__47451;
    wire N__47448;
    wire N__47447;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47431;
    wire N__47430;
    wire N__47427;
    wire N__47426;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47367;
    wire N__47362;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47323;
    wire N__47318;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47303;
    wire N__47296;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47277;
    wire N__47272;
    wire N__47271;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47248;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47224;
    wire N__47221;
    wire N__47216;
    wire N__47213;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__47186;
    wire N__47181;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47171;
    wire N__47166;
    wire N__47163;
    wire N__47158;
    wire N__47155;
    wire N__47154;
    wire N__47151;
    wire N__47148;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47127;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47112;
    wire N__47107;
    wire N__47104;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47094;
    wire N__47089;
    wire N__47088;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47064;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47034;
    wire N__47031;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47014;
    wire N__47011;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46968;
    wire N__46967;
    wire N__46966;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46951;
    wire N__46942;
    wire N__46941;
    wire N__46940;
    wire N__46939;
    wire N__46936;
    wire N__46931;
    wire N__46928;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46912;
    wire N__46911;
    wire N__46908;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46899;
    wire N__46896;
    wire N__46891;
    wire N__46888;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46872;
    wire N__46871;
    wire N__46870;
    wire N__46869;
    wire N__46868;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46862;
    wire N__46853;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46839;
    wire N__46838;
    wire N__46837;
    wire N__46836;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46817;
    wire N__46812;
    wire N__46803;
    wire N__46800;
    wire N__46793;
    wire N__46784;
    wire N__46775;
    wire N__46766;
    wire N__46757;
    wire N__46754;
    wire N__46747;
    wire N__46736;
    wire N__46733;
    wire N__46726;
    wire N__46723;
    wire N__46722;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46699;
    wire N__46696;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46684;
    wire N__46681;
    wire N__46678;
    wire N__46675;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46653;
    wire N__46650;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46633;
    wire N__46630;
    wire N__46627;
    wire N__46626;
    wire N__46625;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46609;
    wire N__46606;
    wire N__46605;
    wire N__46602;
    wire N__46597;
    wire N__46596;
    wire N__46593;
    wire N__46590;
    wire N__46587;
    wire N__46582;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46569;
    wire N__46568;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46552;
    wire N__46549;
    wire N__46548;
    wire N__46547;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46501;
    wire N__46498;
    wire N__46497;
    wire N__46496;
    wire N__46493;
    wire N__46490;
    wire N__46487;
    wire N__46482;
    wire N__46477;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46462;
    wire N__46459;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46447;
    wire N__46444;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46419;
    wire N__46418;
    wire N__46415;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46396;
    wire N__46393;
    wire N__46392;
    wire N__46389;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46359;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46344;
    wire N__46339;
    wire N__46336;
    wire N__46335;
    wire N__46334;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46320;
    wire N__46315;
    wire N__46312;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46300;
    wire N__46297;
    wire N__46296;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46282;
    wire N__46279;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46267;
    wire N__46264;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46249;
    wire N__46246;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46234;
    wire N__46231;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46219;
    wire N__46216;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46204;
    wire N__46201;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46189;
    wire N__46186;
    wire N__46185;
    wire N__46182;
    wire N__46181;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46168;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46147;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46136;
    wire N__46133;
    wire N__46130;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46114;
    wire N__46111;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46099;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46054;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46016;
    wire N__46011;
    wire N__46008;
    wire N__46003;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45961;
    wire N__45958;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45946;
    wire N__45943;
    wire N__45942;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45928;
    wire N__45925;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45908;
    wire N__45901;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45871;
    wire N__45870;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45855;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45840;
    wire N__45837;
    wire N__45836;
    wire N__45835;
    wire N__45834;
    wire N__45833;
    wire N__45832;
    wire N__45829;
    wire N__45828;
    wire N__45827;
    wire N__45826;
    wire N__45825;
    wire N__45824;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45816;
    wire N__45815;
    wire N__45814;
    wire N__45811;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45784;
    wire N__45783;
    wire N__45782;
    wire N__45781;
    wire N__45780;
    wire N__45779;
    wire N__45778;
    wire N__45777;
    wire N__45776;
    wire N__45775;
    wire N__45774;
    wire N__45773;
    wire N__45772;
    wire N__45771;
    wire N__45770;
    wire N__45769;
    wire N__45766;
    wire N__45761;
    wire N__45760;
    wire N__45759;
    wire N__45758;
    wire N__45757;
    wire N__45756;
    wire N__45755;
    wire N__45754;
    wire N__45753;
    wire N__45746;
    wire N__45743;
    wire N__45736;
    wire N__45733;
    wire N__45726;
    wire N__45723;
    wire N__45714;
    wire N__45705;
    wire N__45696;
    wire N__45687;
    wire N__45682;
    wire N__45673;
    wire N__45664;
    wire N__45657;
    wire N__45650;
    wire N__45639;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45606;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45583;
    wire N__45582;
    wire N__45579;
    wire N__45578;
    wire N__45575;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45562;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45541;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45521;
    wire N__45514;
    wire N__45513;
    wire N__45510;
    wire N__45509;
    wire N__45506;
    wire N__45503;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45475;
    wire N__45472;
    wire N__45471;
    wire N__45468;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45451;
    wire N__45450;
    wire N__45447;
    wire N__45446;
    wire N__45443;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45422;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45399;
    wire N__45398;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45378;
    wire N__45373;
    wire N__45370;
    wire N__45369;
    wire N__45366;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45336;
    wire N__45333;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45316;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45300;
    wire N__45297;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45188;
    wire N__45185;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45154;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45130;
    wire N__45129;
    wire N__45128;
    wire N__45125;
    wire N__45120;
    wire N__45115;
    wire N__45112;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44991;
    wire N__44990;
    wire N__44989;
    wire N__44986;
    wire N__44985;
    wire N__44984;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44976;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44968;
    wire N__44961;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44946;
    wire N__44945;
    wire N__44942;
    wire N__44937;
    wire N__44934;
    wire N__44929;
    wire N__44926;
    wire N__44921;
    wire N__44918;
    wire N__44913;
    wire N__44908;
    wire N__44899;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44844;
    wire N__44841;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44804;
    wire N__44799;
    wire N__44796;
    wire N__44795;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44778;
    wire N__44777;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44762;
    wire N__44759;
    wire N__44756;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44740;
    wire N__44739;
    wire N__44736;
    wire N__44735;
    wire N__44734;
    wire N__44733;
    wire N__44730;
    wire N__44729;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44717;
    wire N__44714;
    wire N__44713;
    wire N__44708;
    wire N__44705;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44683;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44671;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44659;
    wire N__44658;
    wire N__44657;
    wire N__44654;
    wire N__44651;
    wire N__44648;
    wire N__44643;
    wire N__44638;
    wire N__44637;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44464;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44419;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44383;
    wire N__44380;
    wire N__44377;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44290;
    wire N__44287;
    wire N__44284;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44216;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44204;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44188;
    wire N__44187;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44177;
    wire N__44172;
    wire N__44167;
    wire N__44164;
    wire N__44163;
    wire N__44160;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44147;
    wire N__44144;
    wire N__44137;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44113;
    wire N__44110;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44091;
    wire N__44088;
    wire N__44087;
    wire N__44084;
    wire N__44081;
    wire N__44078;
    wire N__44071;
    wire N__44070;
    wire N__44069;
    wire N__44066;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44042;
    wire N__44035;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44002;
    wire N__44001;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43914;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43897;
    wire N__43896;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43864;
    wire N__43861;
    wire N__43858;
    wire N__43857;
    wire N__43854;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43825;
    wire N__43822;
    wire N__43821;
    wire N__43818;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43801;
    wire N__43800;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43785;
    wire N__43780;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43772;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43754;
    wire N__43751;
    wire N__43744;
    wire N__43743;
    wire N__43740;
    wire N__43739;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43723;
    wire N__43722;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43707;
    wire N__43706;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43690;
    wire N__43689;
    wire N__43686;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43671;
    wire N__43668;
    wire N__43663;
    wire N__43662;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43643;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43627;
    wire N__43626;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43614;
    wire N__43609;
    wire N__43606;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43598;
    wire N__43597;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43573;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43564;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43506;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43489;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43481;
    wire N__43476;
    wire N__43473;
    wire N__43472;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43453;
    wire N__43450;
    wire N__43449;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43426;
    wire N__43423;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43415;
    wire N__43414;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43398;
    wire N__43395;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43336;
    wire N__43335;
    wire N__43332;
    wire N__43331;
    wire N__43328;
    wire N__43327;
    wire N__43324;
    wire N__43311;
    wire N__43308;
    wire N__43307;
    wire N__43304;
    wire N__43301;
    wire N__43298;
    wire N__43295;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43206;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43189;
    wire N__43188;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42682;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42556;
    wire N__42555;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42505;
    wire N__42502;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42463;
    wire N__42462;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42444;
    wire N__42443;
    wire N__42440;
    wire N__42437;
    wire N__42436;
    wire N__42435;
    wire N__42432;
    wire N__42427;
    wire N__42424;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42412;
    wire N__42409;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42376;
    wire N__42375;
    wire N__42374;
    wire N__42373;
    wire N__42372;
    wire N__42371;
    wire N__42370;
    wire N__42369;
    wire N__42368;
    wire N__42367;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42363;
    wire N__42362;
    wire N__42361;
    wire N__42360;
    wire N__42359;
    wire N__42358;
    wire N__42357;
    wire N__42356;
    wire N__42355;
    wire N__42354;
    wire N__42353;
    wire N__42352;
    wire N__42351;
    wire N__42348;
    wire N__42331;
    wire N__42316;
    wire N__42313;
    wire N__42312;
    wire N__42311;
    wire N__42310;
    wire N__42309;
    wire N__42306;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42291;
    wire N__42284;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42247;
    wire N__42244;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42193;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42181;
    wire N__42180;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42148;
    wire N__42147;
    wire N__42146;
    wire N__42141;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42086;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42074;
    wire N__42067;
    wire N__42064;
    wire N__42061;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42034;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42022;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42009;
    wire N__42006;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41989;
    wire N__41986;
    wire N__41981;
    wire N__41978;
    wire N__41971;
    wire N__41968;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41953;
    wire N__41950;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41902;
    wire N__41899;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41884;
    wire N__41881;
    wire N__41880;
    wire N__41879;
    wire N__41878;
    wire N__41875;
    wire N__41870;
    wire N__41867;
    wire N__41862;
    wire N__41859;
    wire N__41854;
    wire N__41851;
    wire N__41850;
    wire N__41845;
    wire N__41842;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41818;
    wire N__41815;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41803;
    wire N__41802;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41794;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41779;
    wire N__41770;
    wire N__41767;
    wire N__41766;
    wire N__41765;
    wire N__41762;
    wire N__41761;
    wire N__41760;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41734;
    wire N__41731;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41719;
    wire N__41718;
    wire N__41717;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41705;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41680;
    wire N__41679;
    wire N__41678;
    wire N__41673;
    wire N__41670;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41643;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41619;
    wire N__41618;
    wire N__41617;
    wire N__41614;
    wire N__41609;
    wire N__41606;
    wire N__41599;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41587;
    wire N__41584;
    wire N__41583;
    wire N__41582;
    wire N__41579;
    wire N__41578;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41557;
    wire N__41554;
    wire N__41553;
    wire N__41550;
    wire N__41547;
    wire N__41542;
    wire N__41539;
    wire N__41538;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41523;
    wire N__41518;
    wire N__41517;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41494;
    wire N__41493;
    wire N__41490;
    wire N__41489;
    wire N__41486;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41465;
    wire N__41462;
    wire N__41455;
    wire N__41454;
    wire N__41449;
    wire N__41446;
    wire N__41445;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41414;
    wire N__41407;
    wire N__41406;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41383;
    wire N__41380;
    wire N__41379;
    wire N__41374;
    wire N__41371;
    wire N__41370;
    wire N__41365;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41352;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41307;
    wire N__41304;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41296;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41281;
    wire N__41278;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41262;
    wire N__41261;
    wire N__41260;
    wire N__41259;
    wire N__41258;
    wire N__41257;
    wire N__41256;
    wire N__41255;
    wire N__41254;
    wire N__41253;
    wire N__41252;
    wire N__41251;
    wire N__41250;
    wire N__41249;
    wire N__41248;
    wire N__41247;
    wire N__41246;
    wire N__41245;
    wire N__41244;
    wire N__41243;
    wire N__41242;
    wire N__41241;
    wire N__41240;
    wire N__41239;
    wire N__41238;
    wire N__41237;
    wire N__41234;
    wire N__41233;
    wire N__41232;
    wire N__41231;
    wire N__41230;
    wire N__41223;
    wire N__41214;
    wire N__41205;
    wire N__41196;
    wire N__41187;
    wire N__41178;
    wire N__41171;
    wire N__41168;
    wire N__41159;
    wire N__41156;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41067;
    wire N__41062;
    wire N__41059;
    wire N__41058;
    wire N__41055;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41035;
    wire N__41032;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41024;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41008;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40968;
    wire N__40963;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40948;
    wire N__40945;
    wire N__40944;
    wire N__40939;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40924;
    wire N__40921;
    wire N__40920;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40860;
    wire N__40857;
    wire N__40852;
    wire N__40849;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40834;
    wire N__40833;
    wire N__40828;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40800;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40788;
    wire N__40787;
    wire N__40786;
    wire N__40783;
    wire N__40782;
    wire N__40779;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40763;
    wire N__40758;
    wire N__40757;
    wire N__40756;
    wire N__40755;
    wire N__40754;
    wire N__40753;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40744;
    wire N__40741;
    wire N__40740;
    wire N__40737;
    wire N__40736;
    wire N__40733;
    wire N__40732;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40724;
    wire N__40721;
    wire N__40720;
    wire N__40717;
    wire N__40716;
    wire N__40715;
    wire N__40714;
    wire N__40713;
    wire N__40712;
    wire N__40707;
    wire N__40692;
    wire N__40675;
    wire N__40672;
    wire N__40671;
    wire N__40668;
    wire N__40667;
    wire N__40664;
    wire N__40663;
    wire N__40660;
    wire N__40659;
    wire N__40658;
    wire N__40657;
    wire N__40656;
    wire N__40655;
    wire N__40648;
    wire N__40631;
    wire N__40630;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40622;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40613;
    wire N__40612;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40606;
    wire N__40605;
    wire N__40600;
    wire N__40585;
    wire N__40580;
    wire N__40579;
    wire N__40578;
    wire N__40577;
    wire N__40576;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40572;
    wire N__40571;
    wire N__40570;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40556;
    wire N__40547;
    wire N__40546;
    wire N__40539;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40521;
    wire N__40512;
    wire N__40511;
    wire N__40506;
    wire N__40501;
    wire N__40498;
    wire N__40497;
    wire N__40494;
    wire N__40489;
    wire N__40482;
    wire N__40479;
    wire N__40478;
    wire N__40475;
    wire N__40470;
    wire N__40469;
    wire N__40466;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40445;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40427;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40409;
    wire N__40406;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40383;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40366;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40355;
    wire N__40354;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40330;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40216;
    wire N__40213;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40201;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40179;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40131;
    wire N__40126;
    wire N__40123;
    wire N__40120;
    wire N__40117;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40107;
    wire N__40102;
    wire N__40099;
    wire N__40098;
    wire N__40095;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40080;
    wire N__40075;
    wire N__40072;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40060;
    wire N__40057;
    wire N__40056;
    wire N__40051;
    wire N__40048;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40036;
    wire N__40035;
    wire N__40032;
    wire N__40031;
    wire N__40028;
    wire N__40023;
    wire N__40018;
    wire N__40015;
    wire N__40014;
    wire N__40013;
    wire N__40010;
    wire N__40005;
    wire N__40000;
    wire N__39997;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39982;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39916;
    wire N__39915;
    wire N__39912;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39893;
    wire N__39886;
    wire N__39883;
    wire N__39882;
    wire N__39877;
    wire N__39874;
    wire N__39873;
    wire N__39868;
    wire N__39865;
    wire N__39864;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39852;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39829;
    wire N__39828;
    wire N__39823;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39808;
    wire N__39805;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39793;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39771;
    wire N__39766;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39751;
    wire N__39748;
    wire N__39747;
    wire N__39742;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39727;
    wire N__39724;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39713;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39636;
    wire N__39631;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39616;
    wire N__39613;
    wire N__39612;
    wire N__39609;
    wire N__39604;
    wire N__39603;
    wire N__39600;
    wire N__39597;
    wire N__39594;
    wire N__39589;
    wire N__39586;
    wire N__39585;
    wire N__39584;
    wire N__39581;
    wire N__39576;
    wire N__39571;
    wire N__39568;
    wire N__39567;
    wire N__39566;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39550;
    wire N__39547;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39532;
    wire N__39529;
    wire N__39528;
    wire N__39525;
    wire N__39522;
    wire N__39519;
    wire N__39514;
    wire N__39511;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39496;
    wire N__39493;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39478;
    wire N__39475;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39439;
    wire N__39436;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39408;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39382;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39367;
    wire N__39364;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39349;
    wire N__39346;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39331;
    wire N__39328;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39313;
    wire N__39310;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39295;
    wire N__39292;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38937;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38802;
    wire N__38801;
    wire N__38800;
    wire N__38799;
    wire N__38794;
    wire N__38793;
    wire N__38792;
    wire N__38791;
    wire N__38790;
    wire N__38787;
    wire N__38786;
    wire N__38785;
    wire N__38784;
    wire N__38783;
    wire N__38782;
    wire N__38781;
    wire N__38780;
    wire N__38779;
    wire N__38778;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38759;
    wire N__38756;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38738;
    wire N__38737;
    wire N__38736;
    wire N__38735;
    wire N__38734;
    wire N__38733;
    wire N__38732;
    wire N__38731;
    wire N__38730;
    wire N__38729;
    wire N__38728;
    wire N__38721;
    wire N__38712;
    wire N__38709;
    wire N__38708;
    wire N__38703;
    wire N__38700;
    wire N__38699;
    wire N__38694;
    wire N__38683;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38657;
    wire N__38654;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38448;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38417;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38384;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38337;
    wire N__38334;
    wire N__38333;
    wire N__38330;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38257;
    wire N__38254;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38212;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38157;
    wire N__38156;
    wire N__38153;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38040;
    wire N__38037;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38006;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37976;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37952;
    wire N__37947;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37926;
    wire N__37925;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37859;
    wire N__37856;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37823;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37700;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37682;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37656;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37628;
    wire N__37625;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37593;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37560;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37536;
    wire N__37535;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37503;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37483;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37475;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37438;
    wire N__37435;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37383;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37342;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37313;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37267;
    wire N__37264;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37248;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37224;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37190;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37153;
    wire N__37150;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37129;
    wire N__37126;
    wire N__37125;
    wire N__37124;
    wire N__37121;
    wire N__37116;
    wire N__37115;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37050;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37006;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36946;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36915;
    wire N__36914;
    wire N__36911;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36849;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36796;
    wire N__36793;
    wire N__36792;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36780;
    wire N__36775;
    wire N__36772;
    wire N__36771;
    wire N__36768;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36750;
    wire N__36747;
    wire N__36742;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36715;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36685;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36655;
    wire N__36654;
    wire N__36649;
    wire N__36646;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36634;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36582;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36541;
    wire N__36538;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36523;
    wire N__36522;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36505;
    wire N__36502;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36490;
    wire N__36487;
    wire N__36486;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36462;
    wire N__36461;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36399;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36387;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36346;
    wire N__36343;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36333;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36304;
    wire N__36301;
    wire N__36300;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36285;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36273;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36249;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36126;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36102;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36054;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36013;
    wire N__36010;
    wire N__36009;
    wire N__36006;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35989;
    wire N__35988;
    wire N__35985;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35961;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35937;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35913;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35865;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35841;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35787;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35760;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35733;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35718;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35596;
    wire N__35595;
    wire N__35584;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35577;
    wire N__35576;
    wire N__35575;
    wire N__35574;
    wire N__35573;
    wire N__35572;
    wire N__35571;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35566;
    wire N__35565;
    wire N__35564;
    wire N__35563;
    wire N__35562;
    wire N__35557;
    wire N__35554;
    wire N__35553;
    wire N__35552;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35544;
    wire N__35543;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35536;
    wire N__35535;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35520;
    wire N__35513;
    wire N__35502;
    wire N__35501;
    wire N__35500;
    wire N__35499;
    wire N__35498;
    wire N__35497;
    wire N__35496;
    wire N__35493;
    wire N__35486;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35460;
    wire N__35457;
    wire N__35456;
    wire N__35455;
    wire N__35454;
    wire N__35453;
    wire N__35452;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35444;
    wire N__35431;
    wire N__35430;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35423;
    wire N__35422;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35396;
    wire N__35383;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35349;
    wire N__35344;
    wire N__35331;
    wire N__35324;
    wire N__35321;
    wire N__35314;
    wire N__35307;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35245;
    wire N__35244;
    wire N__35243;
    wire N__35242;
    wire N__35241;
    wire N__35240;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35236;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35230;
    wire N__35229;
    wire N__35228;
    wire N__35227;
    wire N__35226;
    wire N__35225;
    wire N__35224;
    wire N__35223;
    wire N__35222;
    wire N__35221;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35215;
    wire N__35210;
    wire N__35199;
    wire N__35198;
    wire N__35197;
    wire N__35194;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35188;
    wire N__35187;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35164;
    wire N__35163;
    wire N__35150;
    wire N__35149;
    wire N__35148;
    wire N__35147;
    wire N__35146;
    wire N__35145;
    wire N__35144;
    wire N__35143;
    wire N__35142;
    wire N__35141;
    wire N__35140;
    wire N__35139;
    wire N__35138;
    wire N__35137;
    wire N__35136;
    wire N__35135;
    wire N__35134;
    wire N__35133;
    wire N__35132;
    wire N__35131;
    wire N__35128;
    wire N__35127;
    wire N__35124;
    wire N__35123;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35115;
    wire N__35114;
    wire N__35113;
    wire N__35112;
    wire N__35111;
    wire N__35110;
    wire N__35109;
    wire N__35108;
    wire N__35093;
    wire N__35088;
    wire N__35085;
    wire N__35080;
    wire N__35077;
    wire N__35076;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35062;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35038;
    wire N__35031;
    wire N__35028;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35016;
    wire N__35015;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35004;
    wire N__35001;
    wire N__35000;
    wire N__34993;
    wire N__34990;
    wire N__34989;
    wire N__34986;
    wire N__34985;
    wire N__34982;
    wire N__34981;
    wire N__34978;
    wire N__34977;
    wire N__34966;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34942;
    wire N__34941;
    wire N__34938;
    wire N__34937;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34929;
    wire N__34926;
    wire N__34925;
    wire N__34922;
    wire N__34921;
    wire N__34918;
    wire N__34911;
    wire N__34908;
    wire N__34903;
    wire N__34902;
    wire N__34901;
    wire N__34900;
    wire N__34897;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34893;
    wire N__34890;
    wire N__34885;
    wire N__34876;
    wire N__34875;
    wire N__34874;
    wire N__34873;
    wire N__34872;
    wire N__34871;
    wire N__34870;
    wire N__34869;
    wire N__34864;
    wire N__34851;
    wire N__34836;
    wire N__34833;
    wire N__34816;
    wire N__34811;
    wire N__34794;
    wire N__34781;
    wire N__34772;
    wire N__34755;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34743;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34735;
    wire N__34732;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34724;
    wire N__34723;
    wire N__34720;
    wire N__34719;
    wire N__34702;
    wire N__34699;
    wire N__34696;
    wire N__34691;
    wire N__34674;
    wire N__34661;
    wire N__34658;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34556;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34479;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34452;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34437;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34384;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34354;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34338;
    wire N__34333;
    wire N__34330;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34303;
    wire N__34300;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34276;
    wire N__34273;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34246;
    wire N__34243;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34210;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34177;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34128;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34098;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34078;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34048;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33994;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33964;
    wire N__33961;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33937;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33904;
    wire N__33903;
    wire N__33900;
    wire N__33895;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33856;
    wire N__33853;
    wire N__33852;
    wire N__33851;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33828;
    wire N__33823;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33808;
    wire N__33805;
    wire N__33804;
    wire N__33803;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33787;
    wire N__33784;
    wire N__33783;
    wire N__33782;
    wire N__33779;
    wire N__33774;
    wire N__33769;
    wire N__33766;
    wire N__33765;
    wire N__33762;
    wire N__33761;
    wire N__33758;
    wire N__33753;
    wire N__33748;
    wire N__33745;
    wire N__33744;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33732;
    wire N__33727;
    wire N__33724;
    wire N__33723;
    wire N__33722;
    wire N__33719;
    wire N__33714;
    wire N__33709;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33682;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33667;
    wire N__33664;
    wire N__33663;
    wire N__33658;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33636;
    wire N__33631;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33609;
    wire N__33604;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33580;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33544;
    wire N__33541;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33529;
    wire N__33526;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33511;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33496;
    wire N__33493;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33481;
    wire N__33478;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33466;
    wire N__33463;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33448;
    wire N__33445;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33430;
    wire N__33427;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33415;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33400;
    wire N__33397;
    wire N__33396;
    wire N__33391;
    wire N__33388;
    wire N__33387;
    wire N__33382;
    wire N__33379;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33306;
    wire N__33305;
    wire N__33304;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33284;
    wire N__33275;
    wire N__33268;
    wire N__33259;
    wire N__33252;
    wire N__33243;
    wire N__33234;
    wire N__33225;
    wire N__33220;
    wire N__33215;
    wire N__33208;
    wire N__33205;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33186;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33143;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33072;
    wire N__33071;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33062;
    wire N__33053;
    wire N__33044;
    wire N__33041;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32970;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32953;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32941;
    wire N__32940;
    wire N__32939;
    wire N__32936;
    wire N__32931;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32881;
    wire N__32880;
    wire N__32879;
    wire N__32878;
    wire N__32877;
    wire N__32876;
    wire N__32875;
    wire N__32874;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32842;
    wire N__32839;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32787;
    wire N__32786;
    wire N__32785;
    wire N__32784;
    wire N__32783;
    wire N__32782;
    wire N__32781;
    wire N__32780;
    wire N__32779;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32764;
    wire N__32763;
    wire N__32762;
    wire N__32761;
    wire N__32748;
    wire N__32745;
    wire N__32744;
    wire N__32743;
    wire N__32740;
    wire N__32735;
    wire N__32728;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32705;
    wire N__32704;
    wire N__32701;
    wire N__32690;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32668;
    wire N__32665;
    wire N__32660;
    wire N__32647;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32635;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32585;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32552;
    wire N__32549;
    wire N__32542;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32534;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32477;
    wire N__32470;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32395;
    wire N__32392;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32377;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32304;
    wire N__32301;
    wire N__32300;
    wire N__32295;
    wire N__32292;
    wire N__32287;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32275;
    wire N__32274;
    wire N__32273;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32160;
    wire N__32155;
    wire N__32152;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32138;
    wire N__32133;
    wire N__32130;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32083;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32056;
    wire N__32053;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32041;
    wire N__32038;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31989;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31965;
    wire N__31960;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31942;
    wire N__31939;
    wire N__31934;
    wire N__31931;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31887;
    wire N__31886;
    wire N__31883;
    wire N__31878;
    wire N__31873;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31865;
    wire N__31862;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31818;
    wire N__31815;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31786;
    wire N__31783;
    wire N__31782;
    wire N__31779;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31761;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31684;
    wire N__31683;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31628;
    wire N__31623;
    wire N__31620;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31603;
    wire N__31600;
    wire N__31599;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31575;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31528;
    wire N__31527;
    wire N__31524;
    wire N__31523;
    wire N__31520;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31508;
    wire N__31503;
    wire N__31500;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31461;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31441;
    wire N__31438;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31425;
    wire N__31422;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31376;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31345;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31287;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31270;
    wire N__31269;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31223;
    wire N__31222;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31142;
    wire N__31141;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31120;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31103;
    wire N__31098;
    wire N__31095;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30976;
    wire N__30973;
    wire N__30972;
    wire N__30971;
    wire N__30968;
    wire N__30963;
    wire N__30958;
    wire N__30957;
    wire N__30952;
    wire N__30949;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30912;
    wire N__30909;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30885;
    wire N__30882;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30821;
    wire N__30814;
    wire N__30813;
    wire N__30810;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30751;
    wire N__30748;
    wire N__30743;
    wire N__30740;
    wire N__30733;
    wire N__30730;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30696;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30669;
    wire N__30668;
    wire N__30665;
    wire N__30660;
    wire N__30659;
    wire N__30654;
    wire N__30651;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30628;
    wire N__30627;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30617;
    wire N__30614;
    wire N__30613;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30585;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30556;
    wire N__30555;
    wire N__30554;
    wire N__30553;
    wire N__30552;
    wire N__30551;
    wire N__30550;
    wire N__30549;
    wire N__30548;
    wire N__30543;
    wire N__30538;
    wire N__30537;
    wire N__30536;
    wire N__30535;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30529;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30523;
    wire N__30516;
    wire N__30505;
    wire N__30504;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30497;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30491;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30467;
    wire N__30462;
    wire N__30455;
    wire N__30442;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30435;
    wire N__30434;
    wire N__30433;
    wire N__30432;
    wire N__30431;
    wire N__30430;
    wire N__30429;
    wire N__30428;
    wire N__30427;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30420;
    wire N__30419;
    wire N__30416;
    wire N__30409;
    wire N__30402;
    wire N__30389;
    wire N__30378;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30358;
    wire N__30357;
    wire N__30356;
    wire N__30347;
    wire N__30346;
    wire N__30343;
    wire N__30336;
    wire N__30331;
    wire N__30330;
    wire N__30329;
    wire N__30328;
    wire N__30327;
    wire N__30326;
    wire N__30325;
    wire N__30324;
    wire N__30323;
    wire N__30322;
    wire N__30321;
    wire N__30320;
    wire N__30319;
    wire N__30306;
    wire N__30305;
    wire N__30304;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30275;
    wire N__30270;
    wire N__30267;
    wire N__30260;
    wire N__30255;
    wire N__30248;
    wire N__30247;
    wire N__30246;
    wire N__30245;
    wire N__30244;
    wire N__30243;
    wire N__30242;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30228;
    wire N__30227;
    wire N__30226;
    wire N__30225;
    wire N__30222;
    wire N__30221;
    wire N__30220;
    wire N__30219;
    wire N__30210;
    wire N__30205;
    wire N__30198;
    wire N__30191;
    wire N__30188;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30172;
    wire N__30165;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30147;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30123;
    wire N__30106;
    wire N__30105;
    wire N__30104;
    wire N__30103;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30099;
    wire N__30098;
    wire N__30097;
    wire N__30096;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30057;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30042;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29953;
    wire N__29950;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29926;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29523;
    wire N__29518;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29494;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29476;
    wire N__29475;
    wire N__29472;
    wire N__29467;
    wire N__29464;
    wire N__29463;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29447;
    wire N__29442;
    wire N__29439;
    wire N__29434;
    wire N__29431;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29419;
    wire N__29418;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29390;
    wire N__29385;
    wire N__29384;
    wire N__29379;
    wire N__29376;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29361;
    wire N__29360;
    wire N__29357;
    wire N__29352;
    wire N__29351;
    wire N__29346;
    wire N__29343;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29265;
    wire N__29260;
    wire N__29257;
    wire N__29256;
    wire N__29255;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29243;
    wire N__29242;
    wire N__29241;
    wire N__29240;
    wire N__29239;
    wire N__29238;
    wire N__29237;
    wire N__29236;
    wire N__29235;
    wire N__29230;
    wire N__29227;
    wire N__29226;
    wire N__29225;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29219;
    wire N__29216;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29196;
    wire N__29195;
    wire N__29194;
    wire N__29193;
    wire N__29192;
    wire N__29191;
    wire N__29190;
    wire N__29189;
    wire N__29188;
    wire N__29187;
    wire N__29186;
    wire N__29183;
    wire N__29174;
    wire N__29167;
    wire N__29164;
    wire N__29159;
    wire N__29150;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29132;
    wire N__29125;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29105;
    wire N__29098;
    wire N__29089;
    wire N__29082;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29063;
    wire N__29058;
    wire N__29055;
    wire N__29046;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29020;
    wire N__28999;
    wire N__28996;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28975;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28951;
    wire N__28948;
    wire N__28947;
    wire N__28946;
    wire N__28945;
    wire N__28942;
    wire N__28935;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28909;
    wire N__28908;
    wire N__28907;
    wire N__28904;
    wire N__28899;
    wire N__28898;
    wire N__28893;
    wire N__28890;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28867;
    wire N__28864;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28819;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28668;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28651;
    wire N__28650;
    wire N__28647;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28609;
    wire N__28606;
    wire N__28605;
    wire N__28604;
    wire N__28603;
    wire N__28600;
    wire N__28595;
    wire N__28592;
    wire N__28585;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28577;
    wire N__28576;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28562;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28383;
    wire N__28382;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28285;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28227;
    wire N__28224;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27474;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27408;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27385;
    wire N__27382;
    wire N__27377;
    wire N__27374;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27322;
    wire N__27319;
    wire N__27314;
    wire N__27311;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27282;
    wire N__27281;
    wire N__27278;
    wire N__27273;
    wire N__27268;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27256;
    wire N__27253;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27241;
    wire N__27240;
    wire N__27235;
    wire N__27232;
    wire N__27231;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27208;
    wire N__27207;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27179;
    wire N__27176;
    wire N__27169;
    wire N__27166;
    wire N__27165;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27152;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27140;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27121;
    wire N__27118;
    wire N__27117;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27097;
    wire N__27096;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27081;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27058;
    wire N__27057;
    wire N__27054;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27019;
    wire N__27016;
    wire N__27015;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27002;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26990;
    wire N__26987;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26971;
    wire N__26968;
    wire N__26967;
    wire N__26964;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26934;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26914;
    wire N__26913;
    wire N__26912;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26880;
    wire N__26875;
    wire N__26874;
    wire N__26869;
    wire N__26866;
    wire N__26865;
    wire N__26862;
    wire N__26861;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26809;
    wire N__26806;
    wire N__26805;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26788;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26743;
    wire N__26742;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26727;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26707;
    wire N__26706;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26686;
    wire N__26683;
    wire N__26678;
    wire N__26675;
    wire N__26668;
    wire N__26665;
    wire N__26664;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26645;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26629;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26617;
    wire N__26616;
    wire N__26615;
    wire N__26612;
    wire N__26607;
    wire N__26602;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26594;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26570;
    wire N__26563;
    wire N__26560;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26539;
    wire N__26538;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26520;
    wire N__26519;
    wire N__26514;
    wire N__26511;
    wire N__26506;
    wire N__26503;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26491;
    wire N__26490;
    wire N__26489;
    wire N__26486;
    wire N__26481;
    wire N__26480;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26461;
    wire N__26460;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26409;
    wire N__26406;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26389;
    wire N__26388;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26350;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26342;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26326;
    wire N__26323;
    wire N__26322;
    wire N__26321;
    wire N__26320;
    wire N__26317;
    wire N__26312;
    wire N__26309;
    wire N__26302;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26287;
    wire N__26286;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26276;
    wire N__26273;
    wire N__26268;
    wire N__26265;
    wire N__26260;
    wire N__26257;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26232;
    wire N__26231;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26215;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26148;
    wire N__26143;
    wire N__26142;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26101;
    wire N__26098;
    wire N__26097;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26085;
    wire N__26080;
    wire N__26077;
    wire N__26076;
    wire N__26073;
    wire N__26072;
    wire N__26069;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26045;
    wire N__26038;
    wire N__26035;
    wire N__26034;
    wire N__26031;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25994;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25953;
    wire N__25952;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25936;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25902;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25890;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25849;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25739;
    wire N__25734;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25629;
    wire N__25624;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25614;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25376;
    wire N__25375;
    wire N__25374;
    wire N__25373;
    wire N__25372;
    wire N__25371;
    wire N__25370;
    wire N__25369;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25362;
    wire N__25361;
    wire N__25360;
    wire N__25359;
    wire N__25358;
    wire N__25357;
    wire N__25356;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25347;
    wire N__25342;
    wire N__25327;
    wire N__25310;
    wire N__25299;
    wire N__25296;
    wire N__25295;
    wire N__25294;
    wire N__25293;
    wire N__25280;
    wire N__25271;
    wire N__25268;
    wire N__25263;
    wire N__25260;
    wire N__25255;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24877;
    wire N__24876;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24856;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24838;
    wire N__24837;
    wire N__24836;
    wire N__24833;
    wire N__24828;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24813;
    wire N__24810;
    wire N__24805;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24729;
    wire N__24726;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24714;
    wire N__24711;
    wire N__24710;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24694;
    wire N__24693;
    wire N__24692;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24663;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24591;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24579;
    wire N__24574;
    wire N__24573;
    wire N__24572;
    wire N__24569;
    wire N__24564;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24091;
    wire N__24090;
    wire N__24087;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24031;
    wire N__24030;
    wire N__24029;
    wire N__24026;
    wire N__24021;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24009;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23992;
    wire N__23989;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23973;
    wire N__23968;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23960;
    wire N__23955;
    wire N__23950;
    wire N__23947;
    wire N__23946;
    wire N__23945;
    wire N__23942;
    wire N__23937;
    wire N__23932;
    wire N__23929;
    wire N__23928;
    wire N__23925;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23902;
    wire N__23899;
    wire N__23898;
    wire N__23895;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23872;
    wire N__23869;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23857;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23836;
    wire N__23833;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23812;
    wire N__23809;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23794;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23770;
    wire N__23767;
    wire N__23766;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23751;
    wire N__23746;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23733;
    wire N__23728;
    wire N__23725;
    wire N__23724;
    wire N__23723;
    wire N__23720;
    wire N__23715;
    wire N__23710;
    wire N__23707;
    wire N__23706;
    wire N__23703;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23680;
    wire N__23677;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23647;
    wire N__23644;
    wire N__23643;
    wire N__23640;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23623;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23604;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23588;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23572;
    wire N__23569;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23548;
    wire N__23545;
    wire N__23544;
    wire N__23541;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23524;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23516;
    wire N__23511;
    wire N__23506;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23498;
    wire N__23493;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23481;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23455;
    wire N__23452;
    wire N__23451;
    wire N__23448;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23241;
    wire N__23236;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23228;
    wire N__23223;
    wire N__23218;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23196;
    wire N__23195;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23108;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23085;
    wire N__23082;
    wire N__23081;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23065;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23028;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23005;
    wire N__23002;
    wire N__23001;
    wire N__23000;
    wire N__22997;
    wire N__22992;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22982;
    wire N__22979;
    wire N__22974;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22923;
    wire N__22922;
    wire N__22921;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22913;
    wire N__22912;
    wire N__22911;
    wire N__22910;
    wire N__22909;
    wire N__22900;
    wire N__22891;
    wire N__22890;
    wire N__22889;
    wire N__22888;
    wire N__22887;
    wire N__22886;
    wire N__22885;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22880;
    wire N__22879;
    wire N__22878;
    wire N__22877;
    wire N__22868;
    wire N__22859;
    wire N__22854;
    wire N__22849;
    wire N__22840;
    wire N__22831;
    wire N__22822;
    wire N__22817;
    wire N__22814;
    wire N__22801;
    wire N__22798;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22762;
    wire N__22761;
    wire N__22760;
    wire N__22757;
    wire N__22756;
    wire N__22753;
    wire N__22748;
    wire N__22745;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22644;
    wire N__22643;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22629;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22573;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22568;
    wire N__22567;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22552;
    wire N__22551;
    wire N__22550;
    wire N__22549;
    wire N__22548;
    wire N__22547;
    wire N__22546;
    wire N__22545;
    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22520;
    wire N__22511;
    wire N__22508;
    wire N__22499;
    wire N__22494;
    wire N__22485;
    wire N__22482;
    wire N__22473;
    wire N__22470;
    wire N__22463;
    wire N__22454;
    wire N__22449;
    wire N__22446;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22410;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22379;
    wire N__22376;
    wire N__22371;
    wire N__22368;
    wire N__22363;
    wire N__22362;
    wire N__22357;
    wire N__22356;
    wire N__22355;
    wire N__22352;
    wire N__22347;
    wire N__22344;
    wire N__22339;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22326;
    wire N__22323;
    wire N__22318;
    wire N__22317;
    wire N__22316;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21976;
    wire N__21973;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21961;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21940;
    wire N__21937;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21925;
    wire N__21924;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21909;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21838;
    wire N__21835;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21784;
    wire N__21781;
    wire N__21780;
    wire N__21779;
    wire N__21776;
    wire N__21771;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21759;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21742;
    wire N__21739;
    wire N__21738;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21723;
    wire N__21718;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21710;
    wire N__21705;
    wire N__21700;
    wire N__21697;
    wire N__21696;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21682;
    wire N__21679;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21652;
    wire N__21649;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21582;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21529;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21521;
    wire N__21516;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21487;
    wire N__21484;
    wire N__21483;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21468;
    wire N__21463;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21450;
    wire N__21445;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21432;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21403;
    wire N__21400;
    wire N__21399;
    wire N__21396;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21371;
    wire N__21366;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21354;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21337;
    wire N__21334;
    wire N__21333;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21318;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21289;
    wire N__21286;
    wire N__21285;
    wire N__21284;
    wire N__21281;
    wire N__21276;
    wire N__21271;
    wire N__21268;
    wire N__21267;
    wire N__21266;
    wire N__21263;
    wire N__21258;
    wire N__21253;
    wire N__21250;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21223;
    wire N__21220;
    wire N__21219;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21145;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21139;
    wire N__21134;
    wire N__21131;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21052;
    wire N__21049;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21034;
    wire N__21031;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21010;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20817;
    wire N__20814;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20778;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20651;
    wire N__20650;
    wire N__20649;
    wire N__20638;
    wire N__20633;
    wire N__20624;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20616;
    wire N__20615;
    wire N__20606;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20594;
    wire N__20583;
    wire N__20580;
    wire N__20575;
    wire N__20572;
    wire N__20563;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20547;
    wire N__20542;
    wire N__20535;
    wire N__20528;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20433;
    wire N__20432;
    wire N__20431;
    wire N__20430;
    wire N__20429;
    wire N__20428;
    wire N__20427;
    wire N__20426;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20421;
    wire N__20420;
    wire N__20419;
    wire N__20418;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20404;
    wire N__20403;
    wire N__20402;
    wire N__20401;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20395;
    wire N__20386;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20378;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20364;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20338;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20313;
    wire N__20304;
    wire N__20299;
    wire N__20286;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19449;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19444;
    wire N__19443;
    wire N__19442;
    wire N__19441;
    wire N__19440;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19393;
    wire N__19384;
    wire N__19379;
    wire N__19374;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire un7_start_stop_0_a3;
    wire bfn_2_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_2_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_2_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_2_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire N_39_i_i;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire bfn_7_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_7_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_7_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_7_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_7_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_7_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire bfn_7_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire bfn_7_17_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.timer_s1.N_161_i ;
    wire delay_hc_input_c_g;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_8_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_8_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_8_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_8_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \delay_measurement_inst.delay_hc_timer.N_199_i ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_198_i ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_8_23_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_8_24_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire bfn_9_7_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_9_8_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_9_9_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_9_10_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.N_1306_i ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_9_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_9_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire s1_phy_c;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_10_8_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_10_9_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire bfn_10_10_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire elapsed_time_ns_1_RNII43T9_0_6_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire bfn_10_14_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_10_15_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_10_16_0_;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_10_17_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_11_20_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_11_21_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire bfn_11_22_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire bfn_11_23_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_11_24_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire bfn_11_25_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire s3_phy_c;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_12_12_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_12_13_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_12_14_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.N_161_i_g ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire bfn_12_26_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_12_27_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire GB_BUFFER_red_c_g_THRU_CO;
    wire bfn_13_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_13_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_13_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_201_i ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire bfn_13_12_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_13_13_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_13_14_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_13_15_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire s2_phy_c;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_13_24_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_13_25_0_;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire bfn_13_26_0_;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire bfn_13_27_0_;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ;
    wire \pwm_generator_inst.threshold_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_14_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_14_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_14_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_14_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_200_i ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire s4_phy_c;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_9_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_15_11_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_15_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_15_14_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_15_15_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire bfn_15_26_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire CONSTANT_ONE_NET;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire bfn_15_27_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_15_28_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.state_RNIE87FZ0Z_2 ;
    wire il_max_comp1_c;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire state_3;
    wire test22_c;
    wire N_19_1;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_16_27_0_;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_16_28_0_;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_16_29_0_;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_17_13_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire test_c;
    wire start_stop_c;
    wire phase_controller_inst1_state_4;
    wire state_ns_i_a3_1;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_17_26_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_17_27_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_17_28_0_;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_18_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_18_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_18_12_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \pwm_generator_inst.N_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \pwm_generator_inst.N_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.N_160 ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire pwm_duty_input_9;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_158 ;
    wire pwm_duty_input_6;
    wire _gnd_net_;
    wire clock_output_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__28675),
            .RESETB(N__33031),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40789),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40577),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__21079,N__34210,N__35644,N__21052,N__21007,N__21193,N__34330,N__29926,N__34177,N__34021,N__34243,N__33960,N__34354,N__34273,N__33937,N__21034}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__40579,dangling_wire_45,N__40578}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40655),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40605),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__42374,N__42367,N__42372,N__42366,N__42373,N__42365,N__42375,N__42362,N__42368,N__42361,N__42369,N__42363,N__42370,N__42364,N__42371}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__40611,N__40608,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__40606,N__40610,N__40607,N__40609}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40576),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40569),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__42351,N__42354,N__42352,N__42355,N__42353,N__50377,N__50323,N__50472,N__50041,N__50266,N__48875,N__48716,N__48958,N__48823,N__50431}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__40575,N__40572,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__40570,N__40574,N__40571,N__40573}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40788),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40782),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__34383,N__34299,N__36684,N__29980,N__36742,N__34407,N__34047,N__31029,N__36714,N__39981,N__34077,N__33993,N__29949,N__46722,N__47880}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__40787,dangling_wire_215,N__40786}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50660),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50662),
            .DIN(N__50661),
            .DOUT(N__50660),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50662),
            .PADOUT(N__50661),
            .PADIN(N__50660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__50651),
            .DIN(N__50650),
            .DOUT(N__50649),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__50651),
            .PADOUT(N__50650),
            .PADIN(N__50649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test_obuf_iopad (
            .OE(N__50642),
            .DIN(N__50641),
            .DOUT(N__50640),
            .PACKAGEPIN(test));
    defparam test_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test_obuf_preio (
            .PADOEN(N__50642),
            .PADOUT(N__50641),
            .PADIN(N__50640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50633),
            .DIN(N__50632),
            .DOUT(N__50631),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50633),
            .PADOUT(N__50632),
            .PADIN(N__50631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50624),
            .DIN(N__50623),
            .DOUT(N__50622),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50624),
            .PADOUT(N__50623),
            .PADIN(N__50622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50615),
            .DIN(N__50614),
            .DOUT(N__50613),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50615),
            .PADOUT(N__50614),
            .PADIN(N__50613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50606),
            .DIN(N__50605),
            .DOUT(N__50604),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50606),
            .PADOUT(N__50605),
            .PADIN(N__50604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50597),
            .DIN(N__50596),
            .DOUT(N__50595),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50597),
            .PADOUT(N__50596),
            .PADIN(N__50595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34144),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test22_obuf_iopad (
            .OE(N__50588),
            .DIN(N__50587),
            .DOUT(N__50586),
            .PACKAGEPIN(test22));
    defparam test22_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test22_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test22_obuf_preio (
            .PADOEN(N__50588),
            .PADOUT(N__50587),
            .PADIN(N__50586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__42400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50579),
            .DIN(N__50578),
            .DOUT(N__50577),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50579),
            .PADOUT(N__50578),
            .PADIN(N__50577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50570),
            .DIN(N__50569),
            .DOUT(N__50568),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50570),
            .PADOUT(N__50569),
            .PADIN(N__50568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50561),
            .DIN(N__50560),
            .DOUT(N__50559),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50561),
            .PADOUT(N__50560),
            .PADIN(N__50559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38920),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50552),
            .DIN(N__50551),
            .DOUT(N__50550),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50552),
            .PADOUT(N__50551),
            .PADIN(N__50550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50543),
            .DIN(N__50542),
            .DOUT(N__50541),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50543),
            .PADOUT(N__50542),
            .PADIN(N__50541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28702),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50534),
            .DIN(N__50533),
            .DOUT(N__50532),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50534),
            .PADOUT(N__50533),
            .PADIN(N__50532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50525),
            .DIN(N__50524),
            .DOUT(N__50523),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50525),
            .PADOUT(N__50524),
            .PADIN(N__50523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__12049 (
            .O(N__50506),
            .I(N__50502));
    InMux I__12048 (
            .O(N__50505),
            .I(N__50498));
    InMux I__12047 (
            .O(N__50502),
            .I(N__50495));
    InMux I__12046 (
            .O(N__50501),
            .I(N__50492));
    LocalMux I__12045 (
            .O(N__50498),
            .I(N__50489));
    LocalMux I__12044 (
            .O(N__50495),
            .I(N__50484));
    LocalMux I__12043 (
            .O(N__50492),
            .I(N__50484));
    Span4Mux_v I__12042 (
            .O(N__50489),
            .I(N__50481));
    Span12Mux_v I__12041 (
            .O(N__50484),
            .I(N__50476));
    Sp12to4 I__12040 (
            .O(N__50481),
            .I(N__50476));
    Odrv12 I__12039 (
            .O(N__50476),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    CascadeMux I__12038 (
            .O(N__50473),
            .I(N__50469));
    InMux I__12037 (
            .O(N__50472),
            .I(N__50465));
    InMux I__12036 (
            .O(N__50469),
            .I(N__50460));
    InMux I__12035 (
            .O(N__50468),
            .I(N__50460));
    LocalMux I__12034 (
            .O(N__50465),
            .I(N__50457));
    LocalMux I__12033 (
            .O(N__50460),
            .I(pwm_duty_input_7));
    Odrv4 I__12032 (
            .O(N__50457),
            .I(pwm_duty_input_7));
    InMux I__12031 (
            .O(N__50452),
            .I(N__50449));
    LocalMux I__12030 (
            .O(N__50449),
            .I(N__50446));
    Odrv4 I__12029 (
            .O(N__50446),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__12028 (
            .O(N__50443),
            .I(N__50434));
    InMux I__12027 (
            .O(N__50442),
            .I(N__50434));
    InMux I__12026 (
            .O(N__50441),
            .I(N__50434));
    LocalMux I__12025 (
            .O(N__50434),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    InMux I__12024 (
            .O(N__50431),
            .I(N__50427));
    InMux I__12023 (
            .O(N__50430),
            .I(N__50424));
    LocalMux I__12022 (
            .O(N__50427),
            .I(N__50421));
    LocalMux I__12021 (
            .O(N__50424),
            .I(pwm_duty_input_0));
    Odrv4 I__12020 (
            .O(N__50421),
            .I(pwm_duty_input_0));
    InMux I__12019 (
            .O(N__50416),
            .I(N__50413));
    LocalMux I__12018 (
            .O(N__50413),
            .I(N__50409));
    InMux I__12017 (
            .O(N__50412),
            .I(N__50406));
    Span4Mux_v I__12016 (
            .O(N__50409),
            .I(N__50400));
    LocalMux I__12015 (
            .O(N__50406),
            .I(N__50400));
    InMux I__12014 (
            .O(N__50405),
            .I(N__50397));
    Span4Mux_v I__12013 (
            .O(N__50400),
            .I(N__50394));
    LocalMux I__12012 (
            .O(N__50397),
            .I(N__50391));
    Sp12to4 I__12011 (
            .O(N__50394),
            .I(N__50388));
    Span4Mux_v I__12010 (
            .O(N__50391),
            .I(N__50385));
    Span12Mux_s3_h I__12009 (
            .O(N__50388),
            .I(N__50380));
    Sp12to4 I__12008 (
            .O(N__50385),
            .I(N__50380));
    Odrv12 I__12007 (
            .O(N__50380),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__12006 (
            .O(N__50377),
            .I(N__50372));
    InMux I__12005 (
            .O(N__50376),
            .I(N__50367));
    InMux I__12004 (
            .O(N__50375),
            .I(N__50367));
    LocalMux I__12003 (
            .O(N__50372),
            .I(N__50364));
    LocalMux I__12002 (
            .O(N__50367),
            .I(pwm_duty_input_9));
    Odrv4 I__12001 (
            .O(N__50364),
            .I(pwm_duty_input_9));
    CascadeMux I__12000 (
            .O(N__50359),
            .I(N__50356));
    InMux I__11999 (
            .O(N__50356),
            .I(N__50353));
    LocalMux I__11998 (
            .O(N__50353),
            .I(N__50349));
    InMux I__11997 (
            .O(N__50352),
            .I(N__50346));
    Span4Mux_v I__11996 (
            .O(N__50349),
            .I(N__50340));
    LocalMux I__11995 (
            .O(N__50346),
            .I(N__50340));
    InMux I__11994 (
            .O(N__50345),
            .I(N__50337));
    Span4Mux_v I__11993 (
            .O(N__50340),
            .I(N__50334));
    LocalMux I__11992 (
            .O(N__50337),
            .I(N__50331));
    Sp12to4 I__11991 (
            .O(N__50334),
            .I(N__50326));
    Span12Mux_v I__11990 (
            .O(N__50331),
            .I(N__50326));
    Odrv12 I__11989 (
            .O(N__50326),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__11988 (
            .O(N__50323),
            .I(N__50318));
    InMux I__11987 (
            .O(N__50322),
            .I(N__50313));
    InMux I__11986 (
            .O(N__50321),
            .I(N__50313));
    LocalMux I__11985 (
            .O(N__50318),
            .I(N__50310));
    LocalMux I__11984 (
            .O(N__50313),
            .I(pwm_duty_input_8));
    Odrv4 I__11983 (
            .O(N__50310),
            .I(pwm_duty_input_8));
    CascadeMux I__11982 (
            .O(N__50305),
            .I(N__50302));
    InMux I__11981 (
            .O(N__50302),
            .I(N__50299));
    LocalMux I__11980 (
            .O(N__50299),
            .I(N__50294));
    InMux I__11979 (
            .O(N__50298),
            .I(N__50291));
    InMux I__11978 (
            .O(N__50297),
            .I(N__50288));
    Span4Mux_v I__11977 (
            .O(N__50294),
            .I(N__50283));
    LocalMux I__11976 (
            .O(N__50291),
            .I(N__50283));
    LocalMux I__11975 (
            .O(N__50288),
            .I(N__50280));
    Span4Mux_v I__11974 (
            .O(N__50283),
            .I(N__50277));
    Span4Mux_v I__11973 (
            .O(N__50280),
            .I(N__50274));
    Sp12to4 I__11972 (
            .O(N__50277),
            .I(N__50269));
    Sp12to4 I__11971 (
            .O(N__50274),
            .I(N__50269));
    Odrv12 I__11970 (
            .O(N__50269),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__11969 (
            .O(N__50266),
            .I(N__50261));
    InMux I__11968 (
            .O(N__50265),
            .I(N__50258));
    InMux I__11967 (
            .O(N__50264),
            .I(N__50255));
    LocalMux I__11966 (
            .O(N__50261),
            .I(N__50252));
    LocalMux I__11965 (
            .O(N__50258),
            .I(pwm_duty_input_5));
    LocalMux I__11964 (
            .O(N__50255),
            .I(pwm_duty_input_5));
    Odrv4 I__11963 (
            .O(N__50252),
            .I(pwm_duty_input_5));
    InMux I__11962 (
            .O(N__50245),
            .I(N__50233));
    InMux I__11961 (
            .O(N__50244),
            .I(N__50230));
    InMux I__11960 (
            .O(N__50243),
            .I(N__50225));
    InMux I__11959 (
            .O(N__50242),
            .I(N__50225));
    InMux I__11958 (
            .O(N__50241),
            .I(N__50222));
    InMux I__11957 (
            .O(N__50240),
            .I(N__50219));
    InMux I__11956 (
            .O(N__50239),
            .I(N__50210));
    InMux I__11955 (
            .O(N__50238),
            .I(N__50210));
    InMux I__11954 (
            .O(N__50237),
            .I(N__50210));
    InMux I__11953 (
            .O(N__50236),
            .I(N__50210));
    LocalMux I__11952 (
            .O(N__50233),
            .I(N__50203));
    LocalMux I__11951 (
            .O(N__50230),
            .I(N__50203));
    LocalMux I__11950 (
            .O(N__50225),
            .I(N__50203));
    LocalMux I__11949 (
            .O(N__50222),
            .I(N__50200));
    LocalMux I__11948 (
            .O(N__50219),
            .I(N__50197));
    LocalMux I__11947 (
            .O(N__50210),
            .I(N__50192));
    Sp12to4 I__11946 (
            .O(N__50203),
            .I(N__50192));
    Span4Mux_h I__11945 (
            .O(N__50200),
            .I(N__50189));
    Span12Mux_s1_h I__11944 (
            .O(N__50197),
            .I(N__50184));
    Span12Mux_s10_v I__11943 (
            .O(N__50192),
            .I(N__50184));
    Odrv4 I__11942 (
            .O(N__50189),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv12 I__11941 (
            .O(N__50184),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__11940 (
            .O(N__50179),
            .I(N__50175));
    InMux I__11939 (
            .O(N__50178),
            .I(N__50171));
    LocalMux I__11938 (
            .O(N__50175),
            .I(N__50168));
    InMux I__11937 (
            .O(N__50174),
            .I(N__50165));
    LocalMux I__11936 (
            .O(N__50171),
            .I(N__50162));
    Span4Mux_v I__11935 (
            .O(N__50168),
            .I(N__50157));
    LocalMux I__11934 (
            .O(N__50165),
            .I(N__50157));
    Span4Mux_v I__11933 (
            .O(N__50162),
            .I(N__50154));
    Span4Mux_v I__11932 (
            .O(N__50157),
            .I(N__50151));
    Sp12to4 I__11931 (
            .O(N__50154),
            .I(N__50146));
    Sp12to4 I__11930 (
            .O(N__50151),
            .I(N__50146));
    Odrv12 I__11929 (
            .O(N__50146),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    CascadeMux I__11928 (
            .O(N__50143),
            .I(N__50137));
    CascadeMux I__11927 (
            .O(N__50142),
            .I(N__50134));
    InMux I__11926 (
            .O(N__50141),
            .I(N__50125));
    InMux I__11925 (
            .O(N__50140),
            .I(N__50125));
    InMux I__11924 (
            .O(N__50137),
            .I(N__50125));
    InMux I__11923 (
            .O(N__50134),
            .I(N__50125));
    LocalMux I__11922 (
            .O(N__50125),
            .I(N__50118));
    InMux I__11921 (
            .O(N__50124),
            .I(N__50115));
    InMux I__11920 (
            .O(N__50123),
            .I(N__50110));
    InMux I__11919 (
            .O(N__50122),
            .I(N__50110));
    InMux I__11918 (
            .O(N__50121),
            .I(N__50107));
    Span4Mux_s2_h I__11917 (
            .O(N__50118),
            .I(N__50100));
    LocalMux I__11916 (
            .O(N__50115),
            .I(N__50100));
    LocalMux I__11915 (
            .O(N__50110),
            .I(N__50100));
    LocalMux I__11914 (
            .O(N__50107),
            .I(N__50097));
    Span4Mux_v I__11913 (
            .O(N__50100),
            .I(N__50094));
    Span12Mux_s10_h I__11912 (
            .O(N__50097),
            .I(N__50091));
    Span4Mux_h I__11911 (
            .O(N__50094),
            .I(N__50088));
    Odrv12 I__11910 (
            .O(N__50091),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__11909 (
            .O(N__50088),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    InMux I__11908 (
            .O(N__50083),
            .I(N__50069));
    InMux I__11907 (
            .O(N__50082),
            .I(N__50069));
    InMux I__11906 (
            .O(N__50081),
            .I(N__50069));
    InMux I__11905 (
            .O(N__50080),
            .I(N__50069));
    InMux I__11904 (
            .O(N__50079),
            .I(N__50064));
    InMux I__11903 (
            .O(N__50078),
            .I(N__50064));
    LocalMux I__11902 (
            .O(N__50069),
            .I(N__50058));
    LocalMux I__11901 (
            .O(N__50064),
            .I(N__50058));
    InMux I__11900 (
            .O(N__50063),
            .I(N__50055));
    Span4Mux_v I__11899 (
            .O(N__50058),
            .I(N__50050));
    LocalMux I__11898 (
            .O(N__50055),
            .I(N__50050));
    Span4Mux_h I__11897 (
            .O(N__50050),
            .I(N__50047));
    Span4Mux_h I__11896 (
            .O(N__50047),
            .I(N__50044));
    Odrv4 I__11895 (
            .O(N__50044),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    InMux I__11894 (
            .O(N__50041),
            .I(N__50036));
    InMux I__11893 (
            .O(N__50040),
            .I(N__50031));
    InMux I__11892 (
            .O(N__50039),
            .I(N__50031));
    LocalMux I__11891 (
            .O(N__50036),
            .I(N__50028));
    LocalMux I__11890 (
            .O(N__50031),
            .I(pwm_duty_input_6));
    Odrv4 I__11889 (
            .O(N__50028),
            .I(pwm_duty_input_6));
    InMux I__11888 (
            .O(N__50023),
            .I(N__50020));
    LocalMux I__11887 (
            .O(N__50020),
            .I(N__49869));
    ClkMux I__11886 (
            .O(N__50019),
            .I(N__49558));
    ClkMux I__11885 (
            .O(N__50018),
            .I(N__49558));
    ClkMux I__11884 (
            .O(N__50017),
            .I(N__49558));
    ClkMux I__11883 (
            .O(N__50016),
            .I(N__49558));
    ClkMux I__11882 (
            .O(N__50015),
            .I(N__49558));
    ClkMux I__11881 (
            .O(N__50014),
            .I(N__49558));
    ClkMux I__11880 (
            .O(N__50013),
            .I(N__49558));
    ClkMux I__11879 (
            .O(N__50012),
            .I(N__49558));
    ClkMux I__11878 (
            .O(N__50011),
            .I(N__49558));
    ClkMux I__11877 (
            .O(N__50010),
            .I(N__49558));
    ClkMux I__11876 (
            .O(N__50009),
            .I(N__49558));
    ClkMux I__11875 (
            .O(N__50008),
            .I(N__49558));
    ClkMux I__11874 (
            .O(N__50007),
            .I(N__49558));
    ClkMux I__11873 (
            .O(N__50006),
            .I(N__49558));
    ClkMux I__11872 (
            .O(N__50005),
            .I(N__49558));
    ClkMux I__11871 (
            .O(N__50004),
            .I(N__49558));
    ClkMux I__11870 (
            .O(N__50003),
            .I(N__49558));
    ClkMux I__11869 (
            .O(N__50002),
            .I(N__49558));
    ClkMux I__11868 (
            .O(N__50001),
            .I(N__49558));
    ClkMux I__11867 (
            .O(N__50000),
            .I(N__49558));
    ClkMux I__11866 (
            .O(N__49999),
            .I(N__49558));
    ClkMux I__11865 (
            .O(N__49998),
            .I(N__49558));
    ClkMux I__11864 (
            .O(N__49997),
            .I(N__49558));
    ClkMux I__11863 (
            .O(N__49996),
            .I(N__49558));
    ClkMux I__11862 (
            .O(N__49995),
            .I(N__49558));
    ClkMux I__11861 (
            .O(N__49994),
            .I(N__49558));
    ClkMux I__11860 (
            .O(N__49993),
            .I(N__49558));
    ClkMux I__11859 (
            .O(N__49992),
            .I(N__49558));
    ClkMux I__11858 (
            .O(N__49991),
            .I(N__49558));
    ClkMux I__11857 (
            .O(N__49990),
            .I(N__49558));
    ClkMux I__11856 (
            .O(N__49989),
            .I(N__49558));
    ClkMux I__11855 (
            .O(N__49988),
            .I(N__49558));
    ClkMux I__11854 (
            .O(N__49987),
            .I(N__49558));
    ClkMux I__11853 (
            .O(N__49986),
            .I(N__49558));
    ClkMux I__11852 (
            .O(N__49985),
            .I(N__49558));
    ClkMux I__11851 (
            .O(N__49984),
            .I(N__49558));
    ClkMux I__11850 (
            .O(N__49983),
            .I(N__49558));
    ClkMux I__11849 (
            .O(N__49982),
            .I(N__49558));
    ClkMux I__11848 (
            .O(N__49981),
            .I(N__49558));
    ClkMux I__11847 (
            .O(N__49980),
            .I(N__49558));
    ClkMux I__11846 (
            .O(N__49979),
            .I(N__49558));
    ClkMux I__11845 (
            .O(N__49978),
            .I(N__49558));
    ClkMux I__11844 (
            .O(N__49977),
            .I(N__49558));
    ClkMux I__11843 (
            .O(N__49976),
            .I(N__49558));
    ClkMux I__11842 (
            .O(N__49975),
            .I(N__49558));
    ClkMux I__11841 (
            .O(N__49974),
            .I(N__49558));
    ClkMux I__11840 (
            .O(N__49973),
            .I(N__49558));
    ClkMux I__11839 (
            .O(N__49972),
            .I(N__49558));
    ClkMux I__11838 (
            .O(N__49971),
            .I(N__49558));
    ClkMux I__11837 (
            .O(N__49970),
            .I(N__49558));
    ClkMux I__11836 (
            .O(N__49969),
            .I(N__49558));
    ClkMux I__11835 (
            .O(N__49968),
            .I(N__49558));
    ClkMux I__11834 (
            .O(N__49967),
            .I(N__49558));
    ClkMux I__11833 (
            .O(N__49966),
            .I(N__49558));
    ClkMux I__11832 (
            .O(N__49965),
            .I(N__49558));
    ClkMux I__11831 (
            .O(N__49964),
            .I(N__49558));
    ClkMux I__11830 (
            .O(N__49963),
            .I(N__49558));
    ClkMux I__11829 (
            .O(N__49962),
            .I(N__49558));
    ClkMux I__11828 (
            .O(N__49961),
            .I(N__49558));
    ClkMux I__11827 (
            .O(N__49960),
            .I(N__49558));
    ClkMux I__11826 (
            .O(N__49959),
            .I(N__49558));
    ClkMux I__11825 (
            .O(N__49958),
            .I(N__49558));
    ClkMux I__11824 (
            .O(N__49957),
            .I(N__49558));
    ClkMux I__11823 (
            .O(N__49956),
            .I(N__49558));
    ClkMux I__11822 (
            .O(N__49955),
            .I(N__49558));
    ClkMux I__11821 (
            .O(N__49954),
            .I(N__49558));
    ClkMux I__11820 (
            .O(N__49953),
            .I(N__49558));
    ClkMux I__11819 (
            .O(N__49952),
            .I(N__49558));
    ClkMux I__11818 (
            .O(N__49951),
            .I(N__49558));
    ClkMux I__11817 (
            .O(N__49950),
            .I(N__49558));
    ClkMux I__11816 (
            .O(N__49949),
            .I(N__49558));
    ClkMux I__11815 (
            .O(N__49948),
            .I(N__49558));
    ClkMux I__11814 (
            .O(N__49947),
            .I(N__49558));
    ClkMux I__11813 (
            .O(N__49946),
            .I(N__49558));
    ClkMux I__11812 (
            .O(N__49945),
            .I(N__49558));
    ClkMux I__11811 (
            .O(N__49944),
            .I(N__49558));
    ClkMux I__11810 (
            .O(N__49943),
            .I(N__49558));
    ClkMux I__11809 (
            .O(N__49942),
            .I(N__49558));
    ClkMux I__11808 (
            .O(N__49941),
            .I(N__49558));
    ClkMux I__11807 (
            .O(N__49940),
            .I(N__49558));
    ClkMux I__11806 (
            .O(N__49939),
            .I(N__49558));
    ClkMux I__11805 (
            .O(N__49938),
            .I(N__49558));
    ClkMux I__11804 (
            .O(N__49937),
            .I(N__49558));
    ClkMux I__11803 (
            .O(N__49936),
            .I(N__49558));
    ClkMux I__11802 (
            .O(N__49935),
            .I(N__49558));
    ClkMux I__11801 (
            .O(N__49934),
            .I(N__49558));
    ClkMux I__11800 (
            .O(N__49933),
            .I(N__49558));
    ClkMux I__11799 (
            .O(N__49932),
            .I(N__49558));
    ClkMux I__11798 (
            .O(N__49931),
            .I(N__49558));
    ClkMux I__11797 (
            .O(N__49930),
            .I(N__49558));
    ClkMux I__11796 (
            .O(N__49929),
            .I(N__49558));
    ClkMux I__11795 (
            .O(N__49928),
            .I(N__49558));
    ClkMux I__11794 (
            .O(N__49927),
            .I(N__49558));
    ClkMux I__11793 (
            .O(N__49926),
            .I(N__49558));
    ClkMux I__11792 (
            .O(N__49925),
            .I(N__49558));
    ClkMux I__11791 (
            .O(N__49924),
            .I(N__49558));
    ClkMux I__11790 (
            .O(N__49923),
            .I(N__49558));
    ClkMux I__11789 (
            .O(N__49922),
            .I(N__49558));
    ClkMux I__11788 (
            .O(N__49921),
            .I(N__49558));
    ClkMux I__11787 (
            .O(N__49920),
            .I(N__49558));
    ClkMux I__11786 (
            .O(N__49919),
            .I(N__49558));
    ClkMux I__11785 (
            .O(N__49918),
            .I(N__49558));
    ClkMux I__11784 (
            .O(N__49917),
            .I(N__49558));
    ClkMux I__11783 (
            .O(N__49916),
            .I(N__49558));
    ClkMux I__11782 (
            .O(N__49915),
            .I(N__49558));
    ClkMux I__11781 (
            .O(N__49914),
            .I(N__49558));
    ClkMux I__11780 (
            .O(N__49913),
            .I(N__49558));
    ClkMux I__11779 (
            .O(N__49912),
            .I(N__49558));
    ClkMux I__11778 (
            .O(N__49911),
            .I(N__49558));
    ClkMux I__11777 (
            .O(N__49910),
            .I(N__49558));
    ClkMux I__11776 (
            .O(N__49909),
            .I(N__49558));
    ClkMux I__11775 (
            .O(N__49908),
            .I(N__49558));
    ClkMux I__11774 (
            .O(N__49907),
            .I(N__49558));
    ClkMux I__11773 (
            .O(N__49906),
            .I(N__49558));
    ClkMux I__11772 (
            .O(N__49905),
            .I(N__49558));
    ClkMux I__11771 (
            .O(N__49904),
            .I(N__49558));
    ClkMux I__11770 (
            .O(N__49903),
            .I(N__49558));
    ClkMux I__11769 (
            .O(N__49902),
            .I(N__49558));
    ClkMux I__11768 (
            .O(N__49901),
            .I(N__49558));
    ClkMux I__11767 (
            .O(N__49900),
            .I(N__49558));
    ClkMux I__11766 (
            .O(N__49899),
            .I(N__49558));
    ClkMux I__11765 (
            .O(N__49898),
            .I(N__49558));
    ClkMux I__11764 (
            .O(N__49897),
            .I(N__49558));
    ClkMux I__11763 (
            .O(N__49896),
            .I(N__49558));
    ClkMux I__11762 (
            .O(N__49895),
            .I(N__49558));
    ClkMux I__11761 (
            .O(N__49894),
            .I(N__49558));
    ClkMux I__11760 (
            .O(N__49893),
            .I(N__49558));
    ClkMux I__11759 (
            .O(N__49892),
            .I(N__49558));
    ClkMux I__11758 (
            .O(N__49891),
            .I(N__49558));
    ClkMux I__11757 (
            .O(N__49890),
            .I(N__49558));
    ClkMux I__11756 (
            .O(N__49889),
            .I(N__49558));
    ClkMux I__11755 (
            .O(N__49888),
            .I(N__49558));
    ClkMux I__11754 (
            .O(N__49887),
            .I(N__49558));
    ClkMux I__11753 (
            .O(N__49886),
            .I(N__49558));
    ClkMux I__11752 (
            .O(N__49885),
            .I(N__49558));
    ClkMux I__11751 (
            .O(N__49884),
            .I(N__49558));
    ClkMux I__11750 (
            .O(N__49883),
            .I(N__49558));
    ClkMux I__11749 (
            .O(N__49882),
            .I(N__49558));
    ClkMux I__11748 (
            .O(N__49881),
            .I(N__49558));
    ClkMux I__11747 (
            .O(N__49880),
            .I(N__49558));
    ClkMux I__11746 (
            .O(N__49879),
            .I(N__49558));
    ClkMux I__11745 (
            .O(N__49878),
            .I(N__49558));
    ClkMux I__11744 (
            .O(N__49877),
            .I(N__49558));
    ClkMux I__11743 (
            .O(N__49876),
            .I(N__49558));
    ClkMux I__11742 (
            .O(N__49875),
            .I(N__49558));
    ClkMux I__11741 (
            .O(N__49874),
            .I(N__49558));
    ClkMux I__11740 (
            .O(N__49873),
            .I(N__49558));
    ClkMux I__11739 (
            .O(N__49872),
            .I(N__49558));
    Glb2LocalMux I__11738 (
            .O(N__49869),
            .I(N__49558));
    ClkMux I__11737 (
            .O(N__49868),
            .I(N__49558));
    ClkMux I__11736 (
            .O(N__49867),
            .I(N__49558));
    ClkMux I__11735 (
            .O(N__49866),
            .I(N__49558));
    ClkMux I__11734 (
            .O(N__49865),
            .I(N__49558));
    GlobalMux I__11733 (
            .O(N__49558),
            .I(clock_output_0));
    InMux I__11732 (
            .O(N__49555),
            .I(N__49549));
    InMux I__11731 (
            .O(N__49554),
            .I(N__49546));
    InMux I__11730 (
            .O(N__49553),
            .I(N__49543));
    InMux I__11729 (
            .O(N__49552),
            .I(N__49540));
    LocalMux I__11728 (
            .O(N__49549),
            .I(N__49537));
    LocalMux I__11727 (
            .O(N__49546),
            .I(N__49534));
    LocalMux I__11726 (
            .O(N__49543),
            .I(N__49531));
    LocalMux I__11725 (
            .O(N__49540),
            .I(N__49527));
    Glb2LocalMux I__11724 (
            .O(N__49537),
            .I(N__49057));
    Glb2LocalMux I__11723 (
            .O(N__49534),
            .I(N__49057));
    Glb2LocalMux I__11722 (
            .O(N__49531),
            .I(N__49057));
    SRMux I__11721 (
            .O(N__49530),
            .I(N__49057));
    Glb2LocalMux I__11720 (
            .O(N__49527),
            .I(N__49057));
    SRMux I__11719 (
            .O(N__49526),
            .I(N__49057));
    SRMux I__11718 (
            .O(N__49525),
            .I(N__49057));
    SRMux I__11717 (
            .O(N__49524),
            .I(N__49057));
    SRMux I__11716 (
            .O(N__49523),
            .I(N__49057));
    SRMux I__11715 (
            .O(N__49522),
            .I(N__49057));
    SRMux I__11714 (
            .O(N__49521),
            .I(N__49057));
    SRMux I__11713 (
            .O(N__49520),
            .I(N__49057));
    SRMux I__11712 (
            .O(N__49519),
            .I(N__49057));
    SRMux I__11711 (
            .O(N__49518),
            .I(N__49057));
    SRMux I__11710 (
            .O(N__49517),
            .I(N__49057));
    SRMux I__11709 (
            .O(N__49516),
            .I(N__49057));
    SRMux I__11708 (
            .O(N__49515),
            .I(N__49057));
    SRMux I__11707 (
            .O(N__49514),
            .I(N__49057));
    SRMux I__11706 (
            .O(N__49513),
            .I(N__49057));
    SRMux I__11705 (
            .O(N__49512),
            .I(N__49057));
    SRMux I__11704 (
            .O(N__49511),
            .I(N__49057));
    SRMux I__11703 (
            .O(N__49510),
            .I(N__49057));
    SRMux I__11702 (
            .O(N__49509),
            .I(N__49057));
    SRMux I__11701 (
            .O(N__49508),
            .I(N__49057));
    SRMux I__11700 (
            .O(N__49507),
            .I(N__49057));
    SRMux I__11699 (
            .O(N__49506),
            .I(N__49057));
    SRMux I__11698 (
            .O(N__49505),
            .I(N__49057));
    SRMux I__11697 (
            .O(N__49504),
            .I(N__49057));
    SRMux I__11696 (
            .O(N__49503),
            .I(N__49057));
    SRMux I__11695 (
            .O(N__49502),
            .I(N__49057));
    SRMux I__11694 (
            .O(N__49501),
            .I(N__49057));
    SRMux I__11693 (
            .O(N__49500),
            .I(N__49057));
    SRMux I__11692 (
            .O(N__49499),
            .I(N__49057));
    SRMux I__11691 (
            .O(N__49498),
            .I(N__49057));
    SRMux I__11690 (
            .O(N__49497),
            .I(N__49057));
    SRMux I__11689 (
            .O(N__49496),
            .I(N__49057));
    SRMux I__11688 (
            .O(N__49495),
            .I(N__49057));
    SRMux I__11687 (
            .O(N__49494),
            .I(N__49057));
    SRMux I__11686 (
            .O(N__49493),
            .I(N__49057));
    SRMux I__11685 (
            .O(N__49492),
            .I(N__49057));
    SRMux I__11684 (
            .O(N__49491),
            .I(N__49057));
    SRMux I__11683 (
            .O(N__49490),
            .I(N__49057));
    SRMux I__11682 (
            .O(N__49489),
            .I(N__49057));
    SRMux I__11681 (
            .O(N__49488),
            .I(N__49057));
    SRMux I__11680 (
            .O(N__49487),
            .I(N__49057));
    SRMux I__11679 (
            .O(N__49486),
            .I(N__49057));
    SRMux I__11678 (
            .O(N__49485),
            .I(N__49057));
    SRMux I__11677 (
            .O(N__49484),
            .I(N__49057));
    SRMux I__11676 (
            .O(N__49483),
            .I(N__49057));
    SRMux I__11675 (
            .O(N__49482),
            .I(N__49057));
    SRMux I__11674 (
            .O(N__49481),
            .I(N__49057));
    SRMux I__11673 (
            .O(N__49480),
            .I(N__49057));
    SRMux I__11672 (
            .O(N__49479),
            .I(N__49057));
    SRMux I__11671 (
            .O(N__49478),
            .I(N__49057));
    SRMux I__11670 (
            .O(N__49477),
            .I(N__49057));
    SRMux I__11669 (
            .O(N__49476),
            .I(N__49057));
    SRMux I__11668 (
            .O(N__49475),
            .I(N__49057));
    SRMux I__11667 (
            .O(N__49474),
            .I(N__49057));
    SRMux I__11666 (
            .O(N__49473),
            .I(N__49057));
    SRMux I__11665 (
            .O(N__49472),
            .I(N__49057));
    SRMux I__11664 (
            .O(N__49471),
            .I(N__49057));
    SRMux I__11663 (
            .O(N__49470),
            .I(N__49057));
    SRMux I__11662 (
            .O(N__49469),
            .I(N__49057));
    SRMux I__11661 (
            .O(N__49468),
            .I(N__49057));
    SRMux I__11660 (
            .O(N__49467),
            .I(N__49057));
    SRMux I__11659 (
            .O(N__49466),
            .I(N__49057));
    SRMux I__11658 (
            .O(N__49465),
            .I(N__49057));
    SRMux I__11657 (
            .O(N__49464),
            .I(N__49057));
    SRMux I__11656 (
            .O(N__49463),
            .I(N__49057));
    SRMux I__11655 (
            .O(N__49462),
            .I(N__49057));
    SRMux I__11654 (
            .O(N__49461),
            .I(N__49057));
    SRMux I__11653 (
            .O(N__49460),
            .I(N__49057));
    SRMux I__11652 (
            .O(N__49459),
            .I(N__49057));
    SRMux I__11651 (
            .O(N__49458),
            .I(N__49057));
    SRMux I__11650 (
            .O(N__49457),
            .I(N__49057));
    SRMux I__11649 (
            .O(N__49456),
            .I(N__49057));
    SRMux I__11648 (
            .O(N__49455),
            .I(N__49057));
    SRMux I__11647 (
            .O(N__49454),
            .I(N__49057));
    SRMux I__11646 (
            .O(N__49453),
            .I(N__49057));
    SRMux I__11645 (
            .O(N__49452),
            .I(N__49057));
    SRMux I__11644 (
            .O(N__49451),
            .I(N__49057));
    SRMux I__11643 (
            .O(N__49450),
            .I(N__49057));
    SRMux I__11642 (
            .O(N__49449),
            .I(N__49057));
    SRMux I__11641 (
            .O(N__49448),
            .I(N__49057));
    SRMux I__11640 (
            .O(N__49447),
            .I(N__49057));
    SRMux I__11639 (
            .O(N__49446),
            .I(N__49057));
    SRMux I__11638 (
            .O(N__49445),
            .I(N__49057));
    SRMux I__11637 (
            .O(N__49444),
            .I(N__49057));
    SRMux I__11636 (
            .O(N__49443),
            .I(N__49057));
    SRMux I__11635 (
            .O(N__49442),
            .I(N__49057));
    SRMux I__11634 (
            .O(N__49441),
            .I(N__49057));
    SRMux I__11633 (
            .O(N__49440),
            .I(N__49057));
    SRMux I__11632 (
            .O(N__49439),
            .I(N__49057));
    SRMux I__11631 (
            .O(N__49438),
            .I(N__49057));
    SRMux I__11630 (
            .O(N__49437),
            .I(N__49057));
    SRMux I__11629 (
            .O(N__49436),
            .I(N__49057));
    SRMux I__11628 (
            .O(N__49435),
            .I(N__49057));
    SRMux I__11627 (
            .O(N__49434),
            .I(N__49057));
    SRMux I__11626 (
            .O(N__49433),
            .I(N__49057));
    SRMux I__11625 (
            .O(N__49432),
            .I(N__49057));
    SRMux I__11624 (
            .O(N__49431),
            .I(N__49057));
    SRMux I__11623 (
            .O(N__49430),
            .I(N__49057));
    SRMux I__11622 (
            .O(N__49429),
            .I(N__49057));
    SRMux I__11621 (
            .O(N__49428),
            .I(N__49057));
    SRMux I__11620 (
            .O(N__49427),
            .I(N__49057));
    SRMux I__11619 (
            .O(N__49426),
            .I(N__49057));
    SRMux I__11618 (
            .O(N__49425),
            .I(N__49057));
    SRMux I__11617 (
            .O(N__49424),
            .I(N__49057));
    SRMux I__11616 (
            .O(N__49423),
            .I(N__49057));
    SRMux I__11615 (
            .O(N__49422),
            .I(N__49057));
    SRMux I__11614 (
            .O(N__49421),
            .I(N__49057));
    SRMux I__11613 (
            .O(N__49420),
            .I(N__49057));
    SRMux I__11612 (
            .O(N__49419),
            .I(N__49057));
    SRMux I__11611 (
            .O(N__49418),
            .I(N__49057));
    SRMux I__11610 (
            .O(N__49417),
            .I(N__49057));
    SRMux I__11609 (
            .O(N__49416),
            .I(N__49057));
    SRMux I__11608 (
            .O(N__49415),
            .I(N__49057));
    SRMux I__11607 (
            .O(N__49414),
            .I(N__49057));
    SRMux I__11606 (
            .O(N__49413),
            .I(N__49057));
    SRMux I__11605 (
            .O(N__49412),
            .I(N__49057));
    SRMux I__11604 (
            .O(N__49411),
            .I(N__49057));
    SRMux I__11603 (
            .O(N__49410),
            .I(N__49057));
    SRMux I__11602 (
            .O(N__49409),
            .I(N__49057));
    SRMux I__11601 (
            .O(N__49408),
            .I(N__49057));
    SRMux I__11600 (
            .O(N__49407),
            .I(N__49057));
    SRMux I__11599 (
            .O(N__49406),
            .I(N__49057));
    SRMux I__11598 (
            .O(N__49405),
            .I(N__49057));
    SRMux I__11597 (
            .O(N__49404),
            .I(N__49057));
    SRMux I__11596 (
            .O(N__49403),
            .I(N__49057));
    SRMux I__11595 (
            .O(N__49402),
            .I(N__49057));
    SRMux I__11594 (
            .O(N__49401),
            .I(N__49057));
    SRMux I__11593 (
            .O(N__49400),
            .I(N__49057));
    SRMux I__11592 (
            .O(N__49399),
            .I(N__49057));
    SRMux I__11591 (
            .O(N__49398),
            .I(N__49057));
    SRMux I__11590 (
            .O(N__49397),
            .I(N__49057));
    SRMux I__11589 (
            .O(N__49396),
            .I(N__49057));
    SRMux I__11588 (
            .O(N__49395),
            .I(N__49057));
    SRMux I__11587 (
            .O(N__49394),
            .I(N__49057));
    SRMux I__11586 (
            .O(N__49393),
            .I(N__49057));
    SRMux I__11585 (
            .O(N__49392),
            .I(N__49057));
    SRMux I__11584 (
            .O(N__49391),
            .I(N__49057));
    SRMux I__11583 (
            .O(N__49390),
            .I(N__49057));
    SRMux I__11582 (
            .O(N__49389),
            .I(N__49057));
    SRMux I__11581 (
            .O(N__49388),
            .I(N__49057));
    SRMux I__11580 (
            .O(N__49387),
            .I(N__49057));
    SRMux I__11579 (
            .O(N__49386),
            .I(N__49057));
    SRMux I__11578 (
            .O(N__49385),
            .I(N__49057));
    SRMux I__11577 (
            .O(N__49384),
            .I(N__49057));
    SRMux I__11576 (
            .O(N__49383),
            .I(N__49057));
    SRMux I__11575 (
            .O(N__49382),
            .I(N__49057));
    SRMux I__11574 (
            .O(N__49381),
            .I(N__49057));
    SRMux I__11573 (
            .O(N__49380),
            .I(N__49057));
    SRMux I__11572 (
            .O(N__49379),
            .I(N__49057));
    SRMux I__11571 (
            .O(N__49378),
            .I(N__49057));
    SRMux I__11570 (
            .O(N__49377),
            .I(N__49057));
    SRMux I__11569 (
            .O(N__49376),
            .I(N__49057));
    SRMux I__11568 (
            .O(N__49375),
            .I(N__49057));
    SRMux I__11567 (
            .O(N__49374),
            .I(N__49057));
    GlobalMux I__11566 (
            .O(N__49057),
            .I(N__49054));
    gio2CtrlBuf I__11565 (
            .O(N__49054),
            .I(red_c_g));
    InMux I__11564 (
            .O(N__49051),
            .I(N__49048));
    LocalMux I__11563 (
            .O(N__49048),
            .I(N__49038));
    InMux I__11562 (
            .O(N__49047),
            .I(N__49023));
    InMux I__11561 (
            .O(N__49046),
            .I(N__49023));
    InMux I__11560 (
            .O(N__49045),
            .I(N__49023));
    InMux I__11559 (
            .O(N__49044),
            .I(N__49023));
    InMux I__11558 (
            .O(N__49043),
            .I(N__49023));
    InMux I__11557 (
            .O(N__49042),
            .I(N__49023));
    InMux I__11556 (
            .O(N__49041),
            .I(N__49023));
    Span4Mux_v I__11555 (
            .O(N__49038),
            .I(N__49018));
    LocalMux I__11554 (
            .O(N__49023),
            .I(N__49018));
    Span4Mux_v I__11553 (
            .O(N__49018),
            .I(N__49013));
    InMux I__11552 (
            .O(N__49017),
            .I(N__49008));
    InMux I__11551 (
            .O(N__49016),
            .I(N__49008));
    Sp12to4 I__11550 (
            .O(N__49013),
            .I(N__49003));
    LocalMux I__11549 (
            .O(N__49008),
            .I(N__49003));
    Span12Mux_h I__11548 (
            .O(N__49003),
            .I(N__49000));
    Odrv12 I__11547 (
            .O(N__49000),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__11546 (
            .O(N__48997),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    InMux I__11545 (
            .O(N__48994),
            .I(N__48991));
    LocalMux I__11544 (
            .O(N__48991),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    CascadeMux I__11543 (
            .O(N__48988),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    CascadeMux I__11542 (
            .O(N__48985),
            .I(N__48982));
    InMux I__11541 (
            .O(N__48982),
            .I(N__48979));
    LocalMux I__11540 (
            .O(N__48979),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__11539 (
            .O(N__48976),
            .I(N__48973));
    LocalMux I__11538 (
            .O(N__48973),
            .I(N__48970));
    Span4Mux_v I__11537 (
            .O(N__48970),
            .I(N__48967));
    Sp12to4 I__11536 (
            .O(N__48967),
            .I(N__48964));
    Span12Mux_s11_h I__11535 (
            .O(N__48964),
            .I(N__48961));
    Odrv12 I__11534 (
            .O(N__48961),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__11533 (
            .O(N__48958),
            .I(N__48955));
    LocalMux I__11532 (
            .O(N__48955),
            .I(N__48951));
    InMux I__11531 (
            .O(N__48954),
            .I(N__48948));
    Span4Mux_v I__11530 (
            .O(N__48951),
            .I(N__48945));
    LocalMux I__11529 (
            .O(N__48948),
            .I(pwm_duty_input_2));
    Odrv4 I__11528 (
            .O(N__48945),
            .I(pwm_duty_input_2));
    InMux I__11527 (
            .O(N__48940),
            .I(N__48937));
    LocalMux I__11526 (
            .O(N__48937),
            .I(N__48934));
    Odrv4 I__11525 (
            .O(N__48934),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__11524 (
            .O(N__48931),
            .I(N__48928));
    LocalMux I__11523 (
            .O(N__48928),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__11522 (
            .O(N__48925),
            .I(N__48920));
    CascadeMux I__11521 (
            .O(N__48924),
            .I(N__48917));
    CascadeMux I__11520 (
            .O(N__48923),
            .I(N__48914));
    InMux I__11519 (
            .O(N__48920),
            .I(N__48911));
    InMux I__11518 (
            .O(N__48917),
            .I(N__48908));
    InMux I__11517 (
            .O(N__48914),
            .I(N__48905));
    LocalMux I__11516 (
            .O(N__48911),
            .I(N__48898));
    LocalMux I__11515 (
            .O(N__48908),
            .I(N__48898));
    LocalMux I__11514 (
            .O(N__48905),
            .I(N__48898));
    Span4Mux_v I__11513 (
            .O(N__48898),
            .I(N__48894));
    InMux I__11512 (
            .O(N__48897),
            .I(N__48891));
    Sp12to4 I__11511 (
            .O(N__48894),
            .I(N__48886));
    LocalMux I__11510 (
            .O(N__48891),
            .I(N__48886));
    Span12Mux_s11_h I__11509 (
            .O(N__48886),
            .I(N__48883));
    Odrv12 I__11508 (
            .O(N__48883),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    CascadeMux I__11507 (
            .O(N__48880),
            .I(N__48877));
    InMux I__11506 (
            .O(N__48877),
            .I(N__48872));
    CascadeMux I__11505 (
            .O(N__48876),
            .I(N__48869));
    InMux I__11504 (
            .O(N__48875),
            .I(N__48866));
    LocalMux I__11503 (
            .O(N__48872),
            .I(N__48863));
    InMux I__11502 (
            .O(N__48869),
            .I(N__48860));
    LocalMux I__11501 (
            .O(N__48866),
            .I(N__48857));
    Span4Mux_h I__11500 (
            .O(N__48863),
            .I(N__48854));
    LocalMux I__11499 (
            .O(N__48860),
            .I(N__48851));
    Span4Mux_v I__11498 (
            .O(N__48857),
            .I(N__48848));
    Odrv4 I__11497 (
            .O(N__48854),
            .I(pwm_duty_input_4));
    Odrv4 I__11496 (
            .O(N__48851),
            .I(pwm_duty_input_4));
    Odrv4 I__11495 (
            .O(N__48848),
            .I(pwm_duty_input_4));
    InMux I__11494 (
            .O(N__48841),
            .I(N__48838));
    LocalMux I__11493 (
            .O(N__48838),
            .I(N__48835));
    Span4Mux_v I__11492 (
            .O(N__48835),
            .I(N__48832));
    Span4Mux_h I__11491 (
            .O(N__48832),
            .I(N__48829));
    Span4Mux_h I__11490 (
            .O(N__48829),
            .I(N__48826));
    Odrv4 I__11489 (
            .O(N__48826),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__11488 (
            .O(N__48823),
            .I(N__48820));
    LocalMux I__11487 (
            .O(N__48820),
            .I(N__48816));
    InMux I__11486 (
            .O(N__48819),
            .I(N__48813));
    Span4Mux_s1_h I__11485 (
            .O(N__48816),
            .I(N__48810));
    LocalMux I__11484 (
            .O(N__48813),
            .I(pwm_duty_input_1));
    Odrv4 I__11483 (
            .O(N__48810),
            .I(pwm_duty_input_1));
    InMux I__11482 (
            .O(N__48805),
            .I(N__48802));
    LocalMux I__11481 (
            .O(N__48802),
            .I(N__48799));
    Span4Mux_v I__11480 (
            .O(N__48799),
            .I(N__48795));
    InMux I__11479 (
            .O(N__48798),
            .I(N__48792));
    Odrv4 I__11478 (
            .O(N__48795),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__11477 (
            .O(N__48792),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__11476 (
            .O(N__48787),
            .I(N__48783));
    InMux I__11475 (
            .O(N__48786),
            .I(N__48780));
    LocalMux I__11474 (
            .O(N__48783),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__11473 (
            .O(N__48780),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__11472 (
            .O(N__48775),
            .I(N__48770));
    InMux I__11471 (
            .O(N__48774),
            .I(N__48767));
    InMux I__11470 (
            .O(N__48773),
            .I(N__48764));
    LocalMux I__11469 (
            .O(N__48770),
            .I(N__48761));
    LocalMux I__11468 (
            .O(N__48767),
            .I(N__48758));
    LocalMux I__11467 (
            .O(N__48764),
            .I(N__48755));
    Span4Mux_v I__11466 (
            .O(N__48761),
            .I(N__48752));
    Span4Mux_s3_h I__11465 (
            .O(N__48758),
            .I(N__48749));
    Span4Mux_s2_h I__11464 (
            .O(N__48755),
            .I(N__48746));
    Sp12to4 I__11463 (
            .O(N__48752),
            .I(N__48743));
    Span4Mux_h I__11462 (
            .O(N__48749),
            .I(N__48740));
    Span4Mux_h I__11461 (
            .O(N__48746),
            .I(N__48737));
    Span12Mux_s11_h I__11460 (
            .O(N__48743),
            .I(N__48734));
    Span4Mux_v I__11459 (
            .O(N__48740),
            .I(N__48731));
    Span4Mux_h I__11458 (
            .O(N__48737),
            .I(N__48728));
    Odrv12 I__11457 (
            .O(N__48734),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__11456 (
            .O(N__48731),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__11455 (
            .O(N__48728),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__11454 (
            .O(N__48721),
            .I(N__48717));
    InMux I__11453 (
            .O(N__48720),
            .I(N__48713));
    LocalMux I__11452 (
            .O(N__48717),
            .I(N__48710));
    InMux I__11451 (
            .O(N__48716),
            .I(N__48707));
    LocalMux I__11450 (
            .O(N__48713),
            .I(N__48704));
    Span4Mux_v I__11449 (
            .O(N__48710),
            .I(N__48701));
    LocalMux I__11448 (
            .O(N__48707),
            .I(N__48698));
    Odrv4 I__11447 (
            .O(N__48704),
            .I(pwm_duty_input_3));
    Odrv4 I__11446 (
            .O(N__48701),
            .I(pwm_duty_input_3));
    Odrv4 I__11445 (
            .O(N__48698),
            .I(pwm_duty_input_3));
    CascadeMux I__11444 (
            .O(N__48691),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__11443 (
            .O(N__48688),
            .I(N__48685));
    LocalMux I__11442 (
            .O(N__48685),
            .I(N__48680));
    InMux I__11441 (
            .O(N__48684),
            .I(N__48675));
    InMux I__11440 (
            .O(N__48683),
            .I(N__48675));
    Odrv4 I__11439 (
            .O(N__48680),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__11438 (
            .O(N__48675),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__11437 (
            .O(N__48670),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__11436 (
            .O(N__48667),
            .I(N__48664));
    LocalMux I__11435 (
            .O(N__48664),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__11434 (
            .O(N__48661),
            .I(N__48658));
    LocalMux I__11433 (
            .O(N__48658),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__11432 (
            .O(N__48655),
            .I(N__48652));
    LocalMux I__11431 (
            .O(N__48652),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__11430 (
            .O(N__48649),
            .I(N__48644));
    InMux I__11429 (
            .O(N__48648),
            .I(N__48641));
    InMux I__11428 (
            .O(N__48647),
            .I(N__48638));
    LocalMux I__11427 (
            .O(N__48644),
            .I(N__48635));
    LocalMux I__11426 (
            .O(N__48641),
            .I(N__48632));
    LocalMux I__11425 (
            .O(N__48638),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv12 I__11424 (
            .O(N__48635),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv4 I__11423 (
            .O(N__48632),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__11422 (
            .O(N__48625),
            .I(N__48620));
    InMux I__11421 (
            .O(N__48624),
            .I(N__48617));
    CascadeMux I__11420 (
            .O(N__48623),
            .I(N__48614));
    LocalMux I__11419 (
            .O(N__48620),
            .I(N__48608));
    LocalMux I__11418 (
            .O(N__48617),
            .I(N__48608));
    InMux I__11417 (
            .O(N__48614),
            .I(N__48605));
    InMux I__11416 (
            .O(N__48613),
            .I(N__48602));
    Span4Mux_v I__11415 (
            .O(N__48608),
            .I(N__48599));
    LocalMux I__11414 (
            .O(N__48605),
            .I(N__48596));
    LocalMux I__11413 (
            .O(N__48602),
            .I(N__48593));
    Span4Mux_h I__11412 (
            .O(N__48599),
            .I(N__48590));
    Span4Mux_v I__11411 (
            .O(N__48596),
            .I(N__48587));
    Odrv4 I__11410 (
            .O(N__48593),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__11409 (
            .O(N__48590),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__11408 (
            .O(N__48587),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__11407 (
            .O(N__48580),
            .I(N__48574));
    InMux I__11406 (
            .O(N__48579),
            .I(N__48574));
    LocalMux I__11405 (
            .O(N__48574),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__11404 (
            .O(N__48571),
            .I(N__48567));
    InMux I__11403 (
            .O(N__48570),
            .I(N__48564));
    InMux I__11402 (
            .O(N__48567),
            .I(N__48561));
    LocalMux I__11401 (
            .O(N__48564),
            .I(N__48558));
    LocalMux I__11400 (
            .O(N__48561),
            .I(N__48555));
    Span4Mux_v I__11399 (
            .O(N__48558),
            .I(N__48551));
    Span4Mux_h I__11398 (
            .O(N__48555),
            .I(N__48548));
    InMux I__11397 (
            .O(N__48554),
            .I(N__48545));
    Span4Mux_h I__11396 (
            .O(N__48551),
            .I(N__48542));
    Span4Mux_h I__11395 (
            .O(N__48548),
            .I(N__48539));
    LocalMux I__11394 (
            .O(N__48545),
            .I(N__48536));
    Span4Mux_h I__11393 (
            .O(N__48542),
            .I(N__48533));
    Span4Mux_h I__11392 (
            .O(N__48539),
            .I(N__48530));
    Span12Mux_h I__11391 (
            .O(N__48536),
            .I(N__48527));
    Span4Mux_v I__11390 (
            .O(N__48533),
            .I(N__48522));
    Span4Mux_v I__11389 (
            .O(N__48530),
            .I(N__48522));
    Odrv12 I__11388 (
            .O(N__48527),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__11387 (
            .O(N__48522),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__11386 (
            .O(N__48517),
            .I(N__48513));
    InMux I__11385 (
            .O(N__48516),
            .I(N__48510));
    LocalMux I__11384 (
            .O(N__48513),
            .I(N__48507));
    LocalMux I__11383 (
            .O(N__48510),
            .I(N__48504));
    Span4Mux_h I__11382 (
            .O(N__48507),
            .I(N__48501));
    Span4Mux_h I__11381 (
            .O(N__48504),
            .I(N__48498));
    Span4Mux_h I__11380 (
            .O(N__48501),
            .I(N__48495));
    Span4Mux_h I__11379 (
            .O(N__48498),
            .I(N__48490));
    Span4Mux_h I__11378 (
            .O(N__48495),
            .I(N__48487));
    InMux I__11377 (
            .O(N__48494),
            .I(N__48482));
    InMux I__11376 (
            .O(N__48493),
            .I(N__48482));
    Span4Mux_h I__11375 (
            .O(N__48490),
            .I(N__48479));
    Span4Mux_v I__11374 (
            .O(N__48487),
            .I(N__48476));
    LocalMux I__11373 (
            .O(N__48482),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__11372 (
            .O(N__48479),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__11371 (
            .O(N__48476),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__11370 (
            .O(N__48469),
            .I(N__48466));
    GlobalMux I__11369 (
            .O(N__48466),
            .I(N__48463));
    gio2CtrlBuf I__11368 (
            .O(N__48463),
            .I(delay_tr_input_c_g));
    InMux I__11367 (
            .O(N__48460),
            .I(N__48455));
    InMux I__11366 (
            .O(N__48459),
            .I(N__48452));
    InMux I__11365 (
            .O(N__48458),
            .I(N__48449));
    LocalMux I__11364 (
            .O(N__48455),
            .I(N__48446));
    LocalMux I__11363 (
            .O(N__48452),
            .I(N__48443));
    LocalMux I__11362 (
            .O(N__48449),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv12 I__11361 (
            .O(N__48446),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv12 I__11360 (
            .O(N__48443),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__11359 (
            .O(N__48436),
            .I(N__48433));
    LocalMux I__11358 (
            .O(N__48433),
            .I(N__48428));
    InMux I__11357 (
            .O(N__48432),
            .I(N__48425));
    InMux I__11356 (
            .O(N__48431),
            .I(N__48422));
    Span4Mux_v I__11355 (
            .O(N__48428),
            .I(N__48414));
    LocalMux I__11354 (
            .O(N__48425),
            .I(N__48414));
    LocalMux I__11353 (
            .O(N__48422),
            .I(N__48414));
    InMux I__11352 (
            .O(N__48421),
            .I(N__48411));
    Span4Mux_h I__11351 (
            .O(N__48414),
            .I(N__48406));
    LocalMux I__11350 (
            .O(N__48411),
            .I(N__48406));
    Span4Mux_h I__11349 (
            .O(N__48406),
            .I(N__48403));
    Odrv4 I__11348 (
            .O(N__48403),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    CascadeMux I__11347 (
            .O(N__48400),
            .I(N__48386));
    InMux I__11346 (
            .O(N__48399),
            .I(N__48375));
    InMux I__11345 (
            .O(N__48398),
            .I(N__48375));
    InMux I__11344 (
            .O(N__48397),
            .I(N__48375));
    InMux I__11343 (
            .O(N__48396),
            .I(N__48366));
    InMux I__11342 (
            .O(N__48395),
            .I(N__48366));
    InMux I__11341 (
            .O(N__48394),
            .I(N__48366));
    InMux I__11340 (
            .O(N__48393),
            .I(N__48366));
    CascadeMux I__11339 (
            .O(N__48392),
            .I(N__48363));
    CascadeMux I__11338 (
            .O(N__48391),
            .I(N__48359));
    InMux I__11337 (
            .O(N__48390),
            .I(N__48339));
    InMux I__11336 (
            .O(N__48389),
            .I(N__48339));
    InMux I__11335 (
            .O(N__48386),
            .I(N__48339));
    InMux I__11334 (
            .O(N__48385),
            .I(N__48339));
    InMux I__11333 (
            .O(N__48384),
            .I(N__48332));
    InMux I__11332 (
            .O(N__48383),
            .I(N__48332));
    InMux I__11331 (
            .O(N__48382),
            .I(N__48332));
    LocalMux I__11330 (
            .O(N__48375),
            .I(N__48310));
    LocalMux I__11329 (
            .O(N__48366),
            .I(N__48310));
    InMux I__11328 (
            .O(N__48363),
            .I(N__48303));
    InMux I__11327 (
            .O(N__48362),
            .I(N__48303));
    InMux I__11326 (
            .O(N__48359),
            .I(N__48303));
    InMux I__11325 (
            .O(N__48358),
            .I(N__48300));
    InMux I__11324 (
            .O(N__48357),
            .I(N__48288));
    InMux I__11323 (
            .O(N__48356),
            .I(N__48288));
    InMux I__11322 (
            .O(N__48355),
            .I(N__48288));
    InMux I__11321 (
            .O(N__48354),
            .I(N__48288));
    InMux I__11320 (
            .O(N__48353),
            .I(N__48285));
    InMux I__11319 (
            .O(N__48352),
            .I(N__48279));
    InMux I__11318 (
            .O(N__48351),
            .I(N__48260));
    InMux I__11317 (
            .O(N__48350),
            .I(N__48260));
    InMux I__11316 (
            .O(N__48349),
            .I(N__48260));
    InMux I__11315 (
            .O(N__48348),
            .I(N__48257));
    LocalMux I__11314 (
            .O(N__48339),
            .I(N__48252));
    LocalMux I__11313 (
            .O(N__48332),
            .I(N__48252));
    InMux I__11312 (
            .O(N__48331),
            .I(N__48247));
    InMux I__11311 (
            .O(N__48330),
            .I(N__48247));
    InMux I__11310 (
            .O(N__48329),
            .I(N__48244));
    InMux I__11309 (
            .O(N__48328),
            .I(N__48239));
    InMux I__11308 (
            .O(N__48327),
            .I(N__48224));
    InMux I__11307 (
            .O(N__48326),
            .I(N__48224));
    InMux I__11306 (
            .O(N__48325),
            .I(N__48224));
    InMux I__11305 (
            .O(N__48324),
            .I(N__48224));
    InMux I__11304 (
            .O(N__48323),
            .I(N__48224));
    InMux I__11303 (
            .O(N__48322),
            .I(N__48224));
    InMux I__11302 (
            .O(N__48321),
            .I(N__48224));
    InMux I__11301 (
            .O(N__48320),
            .I(N__48218));
    InMux I__11300 (
            .O(N__48319),
            .I(N__48215));
    InMux I__11299 (
            .O(N__48318),
            .I(N__48210));
    InMux I__11298 (
            .O(N__48317),
            .I(N__48210));
    InMux I__11297 (
            .O(N__48316),
            .I(N__48207));
    InMux I__11296 (
            .O(N__48315),
            .I(N__48204));
    Span4Mux_h I__11295 (
            .O(N__48310),
            .I(N__48197));
    LocalMux I__11294 (
            .O(N__48303),
            .I(N__48197));
    LocalMux I__11293 (
            .O(N__48300),
            .I(N__48197));
    InMux I__11292 (
            .O(N__48299),
            .I(N__48194));
    InMux I__11291 (
            .O(N__48298),
            .I(N__48191));
    InMux I__11290 (
            .O(N__48297),
            .I(N__48188));
    LocalMux I__11289 (
            .O(N__48288),
            .I(N__48183));
    LocalMux I__11288 (
            .O(N__48285),
            .I(N__48183));
    InMux I__11287 (
            .O(N__48284),
            .I(N__48176));
    InMux I__11286 (
            .O(N__48283),
            .I(N__48176));
    InMux I__11285 (
            .O(N__48282),
            .I(N__48176));
    LocalMux I__11284 (
            .O(N__48279),
            .I(N__48149));
    InMux I__11283 (
            .O(N__48278),
            .I(N__48144));
    InMux I__11282 (
            .O(N__48277),
            .I(N__48144));
    InMux I__11281 (
            .O(N__48276),
            .I(N__48141));
    InMux I__11280 (
            .O(N__48275),
            .I(N__48138));
    InMux I__11279 (
            .O(N__48274),
            .I(N__48135));
    InMux I__11278 (
            .O(N__48273),
            .I(N__48126));
    InMux I__11277 (
            .O(N__48272),
            .I(N__48126));
    InMux I__11276 (
            .O(N__48271),
            .I(N__48126));
    InMux I__11275 (
            .O(N__48270),
            .I(N__48126));
    InMux I__11274 (
            .O(N__48269),
            .I(N__48119));
    InMux I__11273 (
            .O(N__48268),
            .I(N__48119));
    InMux I__11272 (
            .O(N__48267),
            .I(N__48119));
    LocalMux I__11271 (
            .O(N__48260),
            .I(N__48114));
    LocalMux I__11270 (
            .O(N__48257),
            .I(N__48114));
    Span4Mux_h I__11269 (
            .O(N__48252),
            .I(N__48111));
    LocalMux I__11268 (
            .O(N__48247),
            .I(N__48106));
    LocalMux I__11267 (
            .O(N__48244),
            .I(N__48106));
    InMux I__11266 (
            .O(N__48243),
            .I(N__48101));
    InMux I__11265 (
            .O(N__48242),
            .I(N__48101));
    LocalMux I__11264 (
            .O(N__48239),
            .I(N__48096));
    LocalMux I__11263 (
            .O(N__48224),
            .I(N__48096));
    InMux I__11262 (
            .O(N__48223),
            .I(N__48089));
    InMux I__11261 (
            .O(N__48222),
            .I(N__48089));
    InMux I__11260 (
            .O(N__48221),
            .I(N__48089));
    LocalMux I__11259 (
            .O(N__48218),
            .I(N__48084));
    LocalMux I__11258 (
            .O(N__48215),
            .I(N__48084));
    LocalMux I__11257 (
            .O(N__48210),
            .I(N__48081));
    LocalMux I__11256 (
            .O(N__48207),
            .I(N__48078));
    LocalMux I__11255 (
            .O(N__48204),
            .I(N__48075));
    Span4Mux_v I__11254 (
            .O(N__48197),
            .I(N__48072));
    LocalMux I__11253 (
            .O(N__48194),
            .I(N__48061));
    LocalMux I__11252 (
            .O(N__48191),
            .I(N__48061));
    LocalMux I__11251 (
            .O(N__48188),
            .I(N__48061));
    Span4Mux_v I__11250 (
            .O(N__48183),
            .I(N__48061));
    LocalMux I__11249 (
            .O(N__48176),
            .I(N__48061));
    InMux I__11248 (
            .O(N__48175),
            .I(N__48056));
    InMux I__11247 (
            .O(N__48174),
            .I(N__48056));
    InMux I__11246 (
            .O(N__48173),
            .I(N__48049));
    InMux I__11245 (
            .O(N__48172),
            .I(N__48049));
    InMux I__11244 (
            .O(N__48171),
            .I(N__48049));
    InMux I__11243 (
            .O(N__48170),
            .I(N__48044));
    InMux I__11242 (
            .O(N__48169),
            .I(N__48044));
    InMux I__11241 (
            .O(N__48168),
            .I(N__48035));
    InMux I__11240 (
            .O(N__48167),
            .I(N__48035));
    InMux I__11239 (
            .O(N__48166),
            .I(N__48035));
    InMux I__11238 (
            .O(N__48165),
            .I(N__48035));
    InMux I__11237 (
            .O(N__48164),
            .I(N__48032));
    InMux I__11236 (
            .O(N__48163),
            .I(N__48017));
    InMux I__11235 (
            .O(N__48162),
            .I(N__48017));
    InMux I__11234 (
            .O(N__48161),
            .I(N__48017));
    InMux I__11233 (
            .O(N__48160),
            .I(N__48017));
    InMux I__11232 (
            .O(N__48159),
            .I(N__48017));
    InMux I__11231 (
            .O(N__48158),
            .I(N__48017));
    InMux I__11230 (
            .O(N__48157),
            .I(N__48017));
    InMux I__11229 (
            .O(N__48156),
            .I(N__48014));
    InMux I__11228 (
            .O(N__48155),
            .I(N__48007));
    InMux I__11227 (
            .O(N__48154),
            .I(N__48007));
    InMux I__11226 (
            .O(N__48153),
            .I(N__48007));
    InMux I__11225 (
            .O(N__48152),
            .I(N__48004));
    Span4Mux_h I__11224 (
            .O(N__48149),
            .I(N__47999));
    LocalMux I__11223 (
            .O(N__48144),
            .I(N__47999));
    LocalMux I__11222 (
            .O(N__48141),
            .I(N__47996));
    LocalMux I__11221 (
            .O(N__48138),
            .I(N__47985));
    LocalMux I__11220 (
            .O(N__48135),
            .I(N__47985));
    LocalMux I__11219 (
            .O(N__48126),
            .I(N__47985));
    LocalMux I__11218 (
            .O(N__48119),
            .I(N__47985));
    Span4Mux_h I__11217 (
            .O(N__48114),
            .I(N__47985));
    Span4Mux_v I__11216 (
            .O(N__48111),
            .I(N__47980));
    Span4Mux_h I__11215 (
            .O(N__48106),
            .I(N__47980));
    LocalMux I__11214 (
            .O(N__48101),
            .I(N__47961));
    Span4Mux_v I__11213 (
            .O(N__48096),
            .I(N__47961));
    LocalMux I__11212 (
            .O(N__48089),
            .I(N__47961));
    Span4Mux_v I__11211 (
            .O(N__48084),
            .I(N__47961));
    Span4Mux_v I__11210 (
            .O(N__48081),
            .I(N__47961));
    Span4Mux_h I__11209 (
            .O(N__48078),
            .I(N__47961));
    Span4Mux_v I__11208 (
            .O(N__48075),
            .I(N__47961));
    Span4Mux_h I__11207 (
            .O(N__48072),
            .I(N__47961));
    Span4Mux_v I__11206 (
            .O(N__48061),
            .I(N__47961));
    LocalMux I__11205 (
            .O(N__48056),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11204 (
            .O(N__48049),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11203 (
            .O(N__48044),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11202 (
            .O(N__48035),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11201 (
            .O(N__48032),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11200 (
            .O(N__48017),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11199 (
            .O(N__48014),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11198 (
            .O(N__48007),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11197 (
            .O(N__48004),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11196 (
            .O(N__47999),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11195 (
            .O(N__47996),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11194 (
            .O(N__47985),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11193 (
            .O(N__47980),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11192 (
            .O(N__47961),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__11191 (
            .O(N__47932),
            .I(N__47928));
    InMux I__11190 (
            .O(N__47931),
            .I(N__47925));
    LocalMux I__11189 (
            .O(N__47928),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__11188 (
            .O(N__47925),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CEMux I__11187 (
            .O(N__47920),
            .I(N__47890));
    CEMux I__11186 (
            .O(N__47919),
            .I(N__47890));
    CEMux I__11185 (
            .O(N__47918),
            .I(N__47890));
    CEMux I__11184 (
            .O(N__47917),
            .I(N__47890));
    CEMux I__11183 (
            .O(N__47916),
            .I(N__47890));
    CEMux I__11182 (
            .O(N__47915),
            .I(N__47890));
    CEMux I__11181 (
            .O(N__47914),
            .I(N__47890));
    CEMux I__11180 (
            .O(N__47913),
            .I(N__47890));
    CEMux I__11179 (
            .O(N__47912),
            .I(N__47890));
    CEMux I__11178 (
            .O(N__47911),
            .I(N__47890));
    GlobalMux I__11177 (
            .O(N__47890),
            .I(N__47887));
    gio2CtrlBuf I__11176 (
            .O(N__47887),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__11175 (
            .O(N__47884),
            .I(N__47881));
    LocalMux I__11174 (
            .O(N__47881),
            .I(N__47877));
    InMux I__11173 (
            .O(N__47880),
            .I(N__47874));
    Span12Mux_v I__11172 (
            .O(N__47877),
            .I(N__47871));
    LocalMux I__11171 (
            .O(N__47874),
            .I(N__47868));
    Span12Mux_h I__11170 (
            .O(N__47871),
            .I(N__47863));
    Span12Mux_s9_h I__11169 (
            .O(N__47868),
            .I(N__47863));
    Odrv12 I__11168 (
            .O(N__47863),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__11167 (
            .O(N__47860),
            .I(N__47857));
    LocalMux I__11166 (
            .O(N__47857),
            .I(N__47854));
    Span4Mux_v I__11165 (
            .O(N__47854),
            .I(N__47851));
    Odrv4 I__11164 (
            .O(N__47851),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__11163 (
            .O(N__47848),
            .I(N__47845));
    LocalMux I__11162 (
            .O(N__47845),
            .I(N__47835));
    InMux I__11161 (
            .O(N__47844),
            .I(N__47820));
    InMux I__11160 (
            .O(N__47843),
            .I(N__47820));
    InMux I__11159 (
            .O(N__47842),
            .I(N__47820));
    InMux I__11158 (
            .O(N__47841),
            .I(N__47820));
    InMux I__11157 (
            .O(N__47840),
            .I(N__47820));
    InMux I__11156 (
            .O(N__47839),
            .I(N__47820));
    InMux I__11155 (
            .O(N__47838),
            .I(N__47820));
    Span4Mux_v I__11154 (
            .O(N__47835),
            .I(N__47813));
    LocalMux I__11153 (
            .O(N__47820),
            .I(N__47813));
    InMux I__11152 (
            .O(N__47819),
            .I(N__47808));
    InMux I__11151 (
            .O(N__47818),
            .I(N__47808));
    Span4Mux_v I__11150 (
            .O(N__47813),
            .I(N__47803));
    LocalMux I__11149 (
            .O(N__47808),
            .I(N__47803));
    Span4Mux_h I__11148 (
            .O(N__47803),
            .I(N__47800));
    Span4Mux_h I__11147 (
            .O(N__47800),
            .I(N__47797));
    Odrv4 I__11146 (
            .O(N__47797),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__11145 (
            .O(N__47794),
            .I(N__47791));
    InMux I__11144 (
            .O(N__47791),
            .I(N__47788));
    LocalMux I__11143 (
            .O(N__47788),
            .I(N__47785));
    Span4Mux_h I__11142 (
            .O(N__47785),
            .I(N__47782));
    Odrv4 I__11141 (
            .O(N__47782),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    CascadeMux I__11140 (
            .O(N__47779),
            .I(N__47776));
    InMux I__11139 (
            .O(N__47776),
            .I(N__47770));
    InMux I__11138 (
            .O(N__47775),
            .I(N__47770));
    LocalMux I__11137 (
            .O(N__47770),
            .I(N__47766));
    InMux I__11136 (
            .O(N__47769),
            .I(N__47763));
    Span4Mux_h I__11135 (
            .O(N__47766),
            .I(N__47760));
    LocalMux I__11134 (
            .O(N__47763),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__11133 (
            .O(N__47760),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__11132 (
            .O(N__47755),
            .I(N__47750));
    InMux I__11131 (
            .O(N__47754),
            .I(N__47747));
    InMux I__11130 (
            .O(N__47753),
            .I(N__47742));
    InMux I__11129 (
            .O(N__47750),
            .I(N__47742));
    LocalMux I__11128 (
            .O(N__47747),
            .I(N__47737));
    LocalMux I__11127 (
            .O(N__47742),
            .I(N__47737));
    Odrv4 I__11126 (
            .O(N__47737),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__11125 (
            .O(N__47734),
            .I(N__47731));
    LocalMux I__11124 (
            .O(N__47731),
            .I(N__47728));
    Span4Mux_h I__11123 (
            .O(N__47728),
            .I(N__47725));
    Odrv4 I__11122 (
            .O(N__47725),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__11121 (
            .O(N__47722),
            .I(N__47719));
    LocalMux I__11120 (
            .O(N__47719),
            .I(N__47716));
    Span4Mux_h I__11119 (
            .O(N__47716),
            .I(N__47712));
    InMux I__11118 (
            .O(N__47715),
            .I(N__47708));
    Span4Mux_h I__11117 (
            .O(N__47712),
            .I(N__47705));
    InMux I__11116 (
            .O(N__47711),
            .I(N__47702));
    LocalMux I__11115 (
            .O(N__47708),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv4 I__11114 (
            .O(N__47705),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__11113 (
            .O(N__47702),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__11112 (
            .O(N__47695),
            .I(N__47690));
    InMux I__11111 (
            .O(N__47694),
            .I(N__47686));
    CascadeMux I__11110 (
            .O(N__47693),
            .I(N__47683));
    LocalMux I__11109 (
            .O(N__47690),
            .I(N__47680));
    InMux I__11108 (
            .O(N__47689),
            .I(N__47677));
    LocalMux I__11107 (
            .O(N__47686),
            .I(N__47674));
    InMux I__11106 (
            .O(N__47683),
            .I(N__47671));
    Span4Mux_v I__11105 (
            .O(N__47680),
            .I(N__47668));
    LocalMux I__11104 (
            .O(N__47677),
            .I(N__47665));
    Span4Mux_h I__11103 (
            .O(N__47674),
            .I(N__47662));
    LocalMux I__11102 (
            .O(N__47671),
            .I(N__47659));
    Span4Mux_h I__11101 (
            .O(N__47668),
            .I(N__47656));
    Span4Mux_v I__11100 (
            .O(N__47665),
            .I(N__47651));
    Span4Mux_h I__11099 (
            .O(N__47662),
            .I(N__47651));
    Span4Mux_h I__11098 (
            .O(N__47659),
            .I(N__47648));
    Odrv4 I__11097 (
            .O(N__47656),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__11096 (
            .O(N__47651),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__11095 (
            .O(N__47648),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__11094 (
            .O(N__47641),
            .I(N__47635));
    InMux I__11093 (
            .O(N__47640),
            .I(N__47635));
    LocalMux I__11092 (
            .O(N__47635),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__11091 (
            .O(N__47632),
            .I(N__47629));
    LocalMux I__11090 (
            .O(N__47629),
            .I(N__47626));
    Span4Mux_h I__11089 (
            .O(N__47626),
            .I(N__47621));
    InMux I__11088 (
            .O(N__47625),
            .I(N__47618));
    InMux I__11087 (
            .O(N__47624),
            .I(N__47615));
    Span4Mux_h I__11086 (
            .O(N__47621),
            .I(N__47612));
    LocalMux I__11085 (
            .O(N__47618),
            .I(N__47609));
    LocalMux I__11084 (
            .O(N__47615),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__11083 (
            .O(N__47612),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__11082 (
            .O(N__47609),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__11081 (
            .O(N__47602),
            .I(N__47598));
    InMux I__11080 (
            .O(N__47601),
            .I(N__47595));
    LocalMux I__11079 (
            .O(N__47598),
            .I(N__47590));
    LocalMux I__11078 (
            .O(N__47595),
            .I(N__47587));
    InMux I__11077 (
            .O(N__47594),
            .I(N__47584));
    InMux I__11076 (
            .O(N__47593),
            .I(N__47581));
    Span4Mux_h I__11075 (
            .O(N__47590),
            .I(N__47578));
    Span4Mux_h I__11074 (
            .O(N__47587),
            .I(N__47575));
    LocalMux I__11073 (
            .O(N__47584),
            .I(N__47572));
    LocalMux I__11072 (
            .O(N__47581),
            .I(N__47569));
    Span4Mux_v I__11071 (
            .O(N__47578),
            .I(N__47566));
    Span4Mux_h I__11070 (
            .O(N__47575),
            .I(N__47561));
    Span4Mux_v I__11069 (
            .O(N__47572),
            .I(N__47561));
    Odrv12 I__11068 (
            .O(N__47569),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__11067 (
            .O(N__47566),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__11066 (
            .O(N__47561),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__11065 (
            .O(N__47554),
            .I(N__47548));
    InMux I__11064 (
            .O(N__47553),
            .I(N__47548));
    LocalMux I__11063 (
            .O(N__47548),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    InMux I__11062 (
            .O(N__47545),
            .I(N__47540));
    InMux I__11061 (
            .O(N__47544),
            .I(N__47537));
    InMux I__11060 (
            .O(N__47543),
            .I(N__47534));
    LocalMux I__11059 (
            .O(N__47540),
            .I(N__47531));
    LocalMux I__11058 (
            .O(N__47537),
            .I(N__47528));
    LocalMux I__11057 (
            .O(N__47534),
            .I(N__47525));
    Span4Mux_v I__11056 (
            .O(N__47531),
            .I(N__47519));
    Span4Mux_v I__11055 (
            .O(N__47528),
            .I(N__47519));
    Span4Mux_v I__11054 (
            .O(N__47525),
            .I(N__47516));
    InMux I__11053 (
            .O(N__47524),
            .I(N__47513));
    Span4Mux_h I__11052 (
            .O(N__47519),
            .I(N__47510));
    Span4Mux_h I__11051 (
            .O(N__47516),
            .I(N__47507));
    LocalMux I__11050 (
            .O(N__47513),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__11049 (
            .O(N__47510),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__11048 (
            .O(N__47507),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__11047 (
            .O(N__47500),
            .I(N__47497));
    LocalMux I__11046 (
            .O(N__47497),
            .I(N__47493));
    InMux I__11045 (
            .O(N__47496),
            .I(N__47489));
    Span4Mux_h I__11044 (
            .O(N__47493),
            .I(N__47486));
    InMux I__11043 (
            .O(N__47492),
            .I(N__47483));
    LocalMux I__11042 (
            .O(N__47489),
            .I(N__47480));
    Span4Mux_h I__11041 (
            .O(N__47486),
            .I(N__47477));
    LocalMux I__11040 (
            .O(N__47483),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__11039 (
            .O(N__47480),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__11038 (
            .O(N__47477),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__11037 (
            .O(N__47470),
            .I(N__47467));
    LocalMux I__11036 (
            .O(N__47467),
            .I(N__47464));
    Odrv4 I__11035 (
            .O(N__47464),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    InMux I__11034 (
            .O(N__47461),
            .I(N__47455));
    InMux I__11033 (
            .O(N__47460),
            .I(N__47455));
    LocalMux I__11032 (
            .O(N__47455),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    CascadeMux I__11031 (
            .O(N__47452),
            .I(N__47448));
    InMux I__11030 (
            .O(N__47451),
            .I(N__47442));
    InMux I__11029 (
            .O(N__47448),
            .I(N__47442));
    InMux I__11028 (
            .O(N__47447),
            .I(N__47439));
    LocalMux I__11027 (
            .O(N__47442),
            .I(N__47436));
    LocalMux I__11026 (
            .O(N__47439),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__11025 (
            .O(N__47436),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__11024 (
            .O(N__47431),
            .I(N__47427));
    InMux I__11023 (
            .O(N__47430),
            .I(N__47421));
    InMux I__11022 (
            .O(N__47427),
            .I(N__47421));
    InMux I__11021 (
            .O(N__47426),
            .I(N__47418));
    LocalMux I__11020 (
            .O(N__47421),
            .I(N__47415));
    LocalMux I__11019 (
            .O(N__47418),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__11018 (
            .O(N__47415),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    CascadeMux I__11017 (
            .O(N__47410),
            .I(N__47407));
    InMux I__11016 (
            .O(N__47407),
            .I(N__47404));
    LocalMux I__11015 (
            .O(N__47404),
            .I(N__47401));
    Odrv4 I__11014 (
            .O(N__47401),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__11013 (
            .O(N__47398),
            .I(N__47394));
    InMux I__11012 (
            .O(N__47397),
            .I(N__47391));
    LocalMux I__11011 (
            .O(N__47394),
            .I(N__47388));
    LocalMux I__11010 (
            .O(N__47391),
            .I(N__47381));
    Span4Mux_v I__11009 (
            .O(N__47388),
            .I(N__47381));
    InMux I__11008 (
            .O(N__47387),
            .I(N__47378));
    InMux I__11007 (
            .O(N__47386),
            .I(N__47375));
    Span4Mux_h I__11006 (
            .O(N__47381),
            .I(N__47372));
    LocalMux I__11005 (
            .O(N__47378),
            .I(N__47367));
    LocalMux I__11004 (
            .O(N__47375),
            .I(N__47367));
    Odrv4 I__11003 (
            .O(N__47372),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__11002 (
            .O(N__47367),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__11001 (
            .O(N__47362),
            .I(N__47359));
    LocalMux I__11000 (
            .O(N__47359),
            .I(N__47354));
    InMux I__10999 (
            .O(N__47358),
            .I(N__47351));
    InMux I__10998 (
            .O(N__47357),
            .I(N__47348));
    Span4Mux_h I__10997 (
            .O(N__47354),
            .I(N__47345));
    LocalMux I__10996 (
            .O(N__47351),
            .I(N__47342));
    LocalMux I__10995 (
            .O(N__47348),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv4 I__10994 (
            .O(N__47345),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv12 I__10993 (
            .O(N__47342),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__10992 (
            .O(N__47335),
            .I(N__47330));
    InMux I__10991 (
            .O(N__47334),
            .I(N__47327));
    InMux I__10990 (
            .O(N__47333),
            .I(N__47324));
    LocalMux I__10989 (
            .O(N__47330),
            .I(N__47318));
    LocalMux I__10988 (
            .O(N__47327),
            .I(N__47318));
    LocalMux I__10987 (
            .O(N__47324),
            .I(N__47315));
    InMux I__10986 (
            .O(N__47323),
            .I(N__47312));
    Span4Mux_h I__10985 (
            .O(N__47318),
            .I(N__47309));
    Span12Mux_s8_v I__10984 (
            .O(N__47315),
            .I(N__47306));
    LocalMux I__10983 (
            .O(N__47312),
            .I(N__47303));
    Odrv4 I__10982 (
            .O(N__47309),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv12 I__10981 (
            .O(N__47306),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__10980 (
            .O(N__47303),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__10979 (
            .O(N__47296),
            .I(N__47293));
    LocalMux I__10978 (
            .O(N__47293),
            .I(N__47288));
    InMux I__10977 (
            .O(N__47292),
            .I(N__47285));
    InMux I__10976 (
            .O(N__47291),
            .I(N__47282));
    Span4Mux_h I__10975 (
            .O(N__47288),
            .I(N__47277));
    LocalMux I__10974 (
            .O(N__47285),
            .I(N__47277));
    LocalMux I__10973 (
            .O(N__47282),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__10972 (
            .O(N__47277),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__10971 (
            .O(N__47272),
            .I(N__47267));
    InMux I__10970 (
            .O(N__47271),
            .I(N__47264));
    InMux I__10969 (
            .O(N__47270),
            .I(N__47261));
    LocalMux I__10968 (
            .O(N__47267),
            .I(N__47258));
    LocalMux I__10967 (
            .O(N__47264),
            .I(N__47255));
    LocalMux I__10966 (
            .O(N__47261),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__10965 (
            .O(N__47258),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__10964 (
            .O(N__47255),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__10963 (
            .O(N__47248),
            .I(N__47245));
    LocalMux I__10962 (
            .O(N__47245),
            .I(N__47240));
    InMux I__10961 (
            .O(N__47244),
            .I(N__47237));
    InMux I__10960 (
            .O(N__47243),
            .I(N__47234));
    Span4Mux_v I__10959 (
            .O(N__47240),
            .I(N__47231));
    LocalMux I__10958 (
            .O(N__47237),
            .I(N__47228));
    LocalMux I__10957 (
            .O(N__47234),
            .I(N__47225));
    Span4Mux_h I__10956 (
            .O(N__47231),
            .I(N__47221));
    Span4Mux_v I__10955 (
            .O(N__47228),
            .I(N__47216));
    Span4Mux_v I__10954 (
            .O(N__47225),
            .I(N__47216));
    InMux I__10953 (
            .O(N__47224),
            .I(N__47213));
    Odrv4 I__10952 (
            .O(N__47221),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__10951 (
            .O(N__47216),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__10950 (
            .O(N__47213),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__10949 (
            .O(N__47206),
            .I(N__47203));
    LocalMux I__10948 (
            .O(N__47203),
            .I(N__47200));
    Span4Mux_h I__10947 (
            .O(N__47200),
            .I(N__47197));
    Odrv4 I__10946 (
            .O(N__47197),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__10945 (
            .O(N__47194),
            .I(N__47191));
    LocalMux I__10944 (
            .O(N__47191),
            .I(N__47186));
    InMux I__10943 (
            .O(N__47190),
            .I(N__47181));
    InMux I__10942 (
            .O(N__47189),
            .I(N__47181));
    Span4Mux_v I__10941 (
            .O(N__47186),
            .I(N__47177));
    LocalMux I__10940 (
            .O(N__47181),
            .I(N__47174));
    CascadeMux I__10939 (
            .O(N__47180),
            .I(N__47171));
    Span4Mux_h I__10938 (
            .O(N__47177),
            .I(N__47166));
    Span4Mux_v I__10937 (
            .O(N__47174),
            .I(N__47166));
    InMux I__10936 (
            .O(N__47171),
            .I(N__47163));
    Odrv4 I__10935 (
            .O(N__47166),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__10934 (
            .O(N__47163),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__10933 (
            .O(N__47158),
            .I(N__47155));
    LocalMux I__10932 (
            .O(N__47155),
            .I(N__47151));
    InMux I__10931 (
            .O(N__47154),
            .I(N__47148));
    Odrv12 I__10930 (
            .O(N__47151),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__10929 (
            .O(N__47148),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__10928 (
            .O(N__47143),
            .I(N__47140));
    LocalMux I__10927 (
            .O(N__47140),
            .I(N__47137));
    Span4Mux_h I__10926 (
            .O(N__47137),
            .I(N__47134));
    Odrv4 I__10925 (
            .O(N__47134),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__10924 (
            .O(N__47131),
            .I(N__47128));
    InMux I__10923 (
            .O(N__47128),
            .I(N__47123));
    InMux I__10922 (
            .O(N__47127),
            .I(N__47120));
    InMux I__10921 (
            .O(N__47126),
            .I(N__47117));
    LocalMux I__10920 (
            .O(N__47123),
            .I(N__47112));
    LocalMux I__10919 (
            .O(N__47120),
            .I(N__47112));
    LocalMux I__10918 (
            .O(N__47117),
            .I(N__47107));
    Span4Mux_v I__10917 (
            .O(N__47112),
            .I(N__47107));
    Odrv4 I__10916 (
            .O(N__47107),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__10915 (
            .O(N__47104),
            .I(N__47100));
    InMux I__10914 (
            .O(N__47103),
            .I(N__47097));
    LocalMux I__10913 (
            .O(N__47100),
            .I(N__47094));
    LocalMux I__10912 (
            .O(N__47097),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    Odrv4 I__10911 (
            .O(N__47094),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__10910 (
            .O(N__47089),
            .I(N__47085));
    InMux I__10909 (
            .O(N__47088),
            .I(N__47082));
    InMux I__10908 (
            .O(N__47085),
            .I(N__47079));
    LocalMux I__10907 (
            .O(N__47082),
            .I(N__47075));
    LocalMux I__10906 (
            .O(N__47079),
            .I(N__47072));
    InMux I__10905 (
            .O(N__47078),
            .I(N__47069));
    Span4Mux_v I__10904 (
            .O(N__47075),
            .I(N__47064));
    Span4Mux_h I__10903 (
            .O(N__47072),
            .I(N__47064));
    LocalMux I__10902 (
            .O(N__47069),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__10901 (
            .O(N__47064),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__10900 (
            .O(N__47059),
            .I(N__47056));
    InMux I__10899 (
            .O(N__47056),
            .I(N__47053));
    LocalMux I__10898 (
            .O(N__47053),
            .I(N__47050));
    Span4Mux_h I__10897 (
            .O(N__47050),
            .I(N__47047));
    Span4Mux_h I__10896 (
            .O(N__47047),
            .I(N__47044));
    Odrv4 I__10895 (
            .O(N__47044),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__10894 (
            .O(N__47041),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__10893 (
            .O(N__47038),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__10892 (
            .O(N__47035),
            .I(N__47031));
    InMux I__10891 (
            .O(N__47034),
            .I(N__47027));
    LocalMux I__10890 (
            .O(N__47031),
            .I(N__47024));
    InMux I__10889 (
            .O(N__47030),
            .I(N__47021));
    LocalMux I__10888 (
            .O(N__47027),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__10887 (
            .O(N__47024),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    LocalMux I__10886 (
            .O(N__47021),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__10885 (
            .O(N__47014),
            .I(N__47011));
    LocalMux I__10884 (
            .O(N__47011),
            .I(N__47007));
    InMux I__10883 (
            .O(N__47010),
            .I(N__47004));
    Odrv4 I__10882 (
            .O(N__47007),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__10881 (
            .O(N__47004),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__10880 (
            .O(N__46999),
            .I(N__46996));
    InMux I__10879 (
            .O(N__46996),
            .I(N__46993));
    LocalMux I__10878 (
            .O(N__46993),
            .I(N__46990));
    Odrv12 I__10877 (
            .O(N__46990),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__10876 (
            .O(N__46987),
            .I(N__46983));
    InMux I__10875 (
            .O(N__46986),
            .I(N__46980));
    LocalMux I__10874 (
            .O(N__46983),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__10873 (
            .O(N__46980),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__10872 (
            .O(N__46975),
            .I(N__46972));
    LocalMux I__10871 (
            .O(N__46972),
            .I(N__46969));
    Span4Mux_h I__10870 (
            .O(N__46969),
            .I(N__46962));
    InMux I__10869 (
            .O(N__46968),
            .I(N__46959));
    InMux I__10868 (
            .O(N__46967),
            .I(N__46956));
    InMux I__10867 (
            .O(N__46966),
            .I(N__46951));
    InMux I__10866 (
            .O(N__46965),
            .I(N__46951));
    Odrv4 I__10865 (
            .O(N__46962),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__10864 (
            .O(N__46959),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__10863 (
            .O(N__46956),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__10862 (
            .O(N__46951),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__10861 (
            .O(N__46942),
            .I(N__46936));
    InMux I__10860 (
            .O(N__46941),
            .I(N__46931));
    InMux I__10859 (
            .O(N__46940),
            .I(N__46931));
    CascadeMux I__10858 (
            .O(N__46939),
            .I(N__46928));
    LocalMux I__10857 (
            .O(N__46936),
            .I(N__46923));
    LocalMux I__10856 (
            .O(N__46931),
            .I(N__46923));
    InMux I__10855 (
            .O(N__46928),
            .I(N__46920));
    Span4Mux_v I__10854 (
            .O(N__46923),
            .I(N__46917));
    LocalMux I__10853 (
            .O(N__46920),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__10852 (
            .O(N__46917),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__10851 (
            .O(N__46912),
            .I(N__46908));
    CascadeMux I__10850 (
            .O(N__46911),
            .I(N__46905));
    InMux I__10849 (
            .O(N__46908),
            .I(N__46899));
    InMux I__10848 (
            .O(N__46905),
            .I(N__46896));
    InMux I__10847 (
            .O(N__46904),
            .I(N__46891));
    InMux I__10846 (
            .O(N__46903),
            .I(N__46891));
    InMux I__10845 (
            .O(N__46902),
            .I(N__46888));
    LocalMux I__10844 (
            .O(N__46899),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__10843 (
            .O(N__46896),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__10842 (
            .O(N__46891),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__10841 (
            .O(N__46888),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    IoInMux I__10840 (
            .O(N__46879),
            .I(N__46876));
    LocalMux I__10839 (
            .O(N__46876),
            .I(N__46873));
    IoSpan4Mux I__10838 (
            .O(N__46873),
            .I(N__46862));
    InMux I__10837 (
            .O(N__46872),
            .I(N__46853));
    InMux I__10836 (
            .O(N__46871),
            .I(N__46853));
    InMux I__10835 (
            .O(N__46870),
            .I(N__46853));
    InMux I__10834 (
            .O(N__46869),
            .I(N__46853));
    InMux I__10833 (
            .O(N__46868),
            .I(N__46846));
    InMux I__10832 (
            .O(N__46867),
            .I(N__46846));
    InMux I__10831 (
            .O(N__46866),
            .I(N__46846));
    InMux I__10830 (
            .O(N__46865),
            .I(N__46839));
    Span4Mux_s3_v I__10829 (
            .O(N__46862),
            .I(N__46817));
    LocalMux I__10828 (
            .O(N__46853),
            .I(N__46812));
    LocalMux I__10827 (
            .O(N__46846),
            .I(N__46812));
    InMux I__10826 (
            .O(N__46845),
            .I(N__46803));
    InMux I__10825 (
            .O(N__46844),
            .I(N__46803));
    InMux I__10824 (
            .O(N__46843),
            .I(N__46803));
    InMux I__10823 (
            .O(N__46842),
            .I(N__46803));
    LocalMux I__10822 (
            .O(N__46839),
            .I(N__46800));
    InMux I__10821 (
            .O(N__46838),
            .I(N__46793));
    InMux I__10820 (
            .O(N__46837),
            .I(N__46793));
    InMux I__10819 (
            .O(N__46836),
            .I(N__46793));
    InMux I__10818 (
            .O(N__46835),
            .I(N__46784));
    InMux I__10817 (
            .O(N__46834),
            .I(N__46784));
    InMux I__10816 (
            .O(N__46833),
            .I(N__46784));
    InMux I__10815 (
            .O(N__46832),
            .I(N__46784));
    InMux I__10814 (
            .O(N__46831),
            .I(N__46775));
    InMux I__10813 (
            .O(N__46830),
            .I(N__46775));
    InMux I__10812 (
            .O(N__46829),
            .I(N__46775));
    InMux I__10811 (
            .O(N__46828),
            .I(N__46775));
    InMux I__10810 (
            .O(N__46827),
            .I(N__46766));
    InMux I__10809 (
            .O(N__46826),
            .I(N__46766));
    InMux I__10808 (
            .O(N__46825),
            .I(N__46766));
    InMux I__10807 (
            .O(N__46824),
            .I(N__46766));
    InMux I__10806 (
            .O(N__46823),
            .I(N__46757));
    InMux I__10805 (
            .O(N__46822),
            .I(N__46757));
    InMux I__10804 (
            .O(N__46821),
            .I(N__46757));
    InMux I__10803 (
            .O(N__46820),
            .I(N__46757));
    Sp12to4 I__10802 (
            .O(N__46817),
            .I(N__46754));
    Span4Mux_v I__10801 (
            .O(N__46812),
            .I(N__46747));
    LocalMux I__10800 (
            .O(N__46803),
            .I(N__46747));
    Span4Mux_h I__10799 (
            .O(N__46800),
            .I(N__46747));
    LocalMux I__10798 (
            .O(N__46793),
            .I(N__46736));
    LocalMux I__10797 (
            .O(N__46784),
            .I(N__46736));
    LocalMux I__10796 (
            .O(N__46775),
            .I(N__46736));
    LocalMux I__10795 (
            .O(N__46766),
            .I(N__46736));
    LocalMux I__10794 (
            .O(N__46757),
            .I(N__46736));
    Span12Mux_v I__10793 (
            .O(N__46754),
            .I(N__46733));
    Odrv4 I__10792 (
            .O(N__46747),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__10791 (
            .O(N__46736),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__10790 (
            .O(N__46733),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__10789 (
            .O(N__46726),
            .I(N__46723));
    LocalMux I__10788 (
            .O(N__46723),
            .I(N__46719));
    InMux I__10787 (
            .O(N__46722),
            .I(N__46716));
    Span4Mux_h I__10786 (
            .O(N__46719),
            .I(N__46713));
    LocalMux I__10785 (
            .O(N__46716),
            .I(N__46710));
    Span4Mux_h I__10784 (
            .O(N__46713),
            .I(N__46707));
    Span4Mux_s3_h I__10783 (
            .O(N__46710),
            .I(N__46704));
    Span4Mux_h I__10782 (
            .O(N__46707),
            .I(N__46699));
    Span4Mux_h I__10781 (
            .O(N__46704),
            .I(N__46699));
    Odrv4 I__10780 (
            .O(N__46699),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__10779 (
            .O(N__46696),
            .I(N__46692));
    InMux I__10778 (
            .O(N__46695),
            .I(N__46689));
    LocalMux I__10777 (
            .O(N__46692),
            .I(N__46684));
    LocalMux I__10776 (
            .O(N__46689),
            .I(N__46684));
    Span4Mux_v I__10775 (
            .O(N__46684),
            .I(N__46681));
    Odrv4 I__10774 (
            .O(N__46681),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__10773 (
            .O(N__46678),
            .I(N__46675));
    LocalMux I__10772 (
            .O(N__46675),
            .I(N__46671));
    InMux I__10771 (
            .O(N__46674),
            .I(N__46668));
    Span4Mux_h I__10770 (
            .O(N__46671),
            .I(N__46663));
    LocalMux I__10769 (
            .O(N__46668),
            .I(N__46663));
    Span4Mux_h I__10768 (
            .O(N__46663),
            .I(N__46660));
    Span4Mux_h I__10767 (
            .O(N__46660),
            .I(N__46657));
    Odrv4 I__10766 (
            .O(N__46657),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__10765 (
            .O(N__46654),
            .I(N__46650));
    InMux I__10764 (
            .O(N__46653),
            .I(N__46646));
    LocalMux I__10763 (
            .O(N__46650),
            .I(N__46643));
    InMux I__10762 (
            .O(N__46649),
            .I(N__46640));
    LocalMux I__10761 (
            .O(N__46646),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv12 I__10760 (
            .O(N__46643),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    LocalMux I__10759 (
            .O(N__46640),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    IoInMux I__10758 (
            .O(N__46633),
            .I(N__46630));
    LocalMux I__10757 (
            .O(N__46630),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__10756 (
            .O(N__46627),
            .I(N__46620));
    InMux I__10755 (
            .O(N__46626),
            .I(N__46620));
    InMux I__10754 (
            .O(N__46625),
            .I(N__46617));
    LocalMux I__10753 (
            .O(N__46620),
            .I(N__46614));
    LocalMux I__10752 (
            .O(N__46617),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__10751 (
            .O(N__46614),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__10750 (
            .O(N__46609),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    CascadeMux I__10749 (
            .O(N__46606),
            .I(N__46602));
    InMux I__10748 (
            .O(N__46605),
            .I(N__46597));
    InMux I__10747 (
            .O(N__46602),
            .I(N__46597));
    LocalMux I__10746 (
            .O(N__46597),
            .I(N__46593));
    InMux I__10745 (
            .O(N__46596),
            .I(N__46590));
    Span4Mux_h I__10744 (
            .O(N__46593),
            .I(N__46587));
    LocalMux I__10743 (
            .O(N__46590),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__10742 (
            .O(N__46587),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__10741 (
            .O(N__46582),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__10740 (
            .O(N__46579),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__10739 (
            .O(N__46576),
            .I(bfn_18_13_0_));
    CascadeMux I__10738 (
            .O(N__46573),
            .I(N__46570));
    InMux I__10737 (
            .O(N__46570),
            .I(N__46563));
    InMux I__10736 (
            .O(N__46569),
            .I(N__46563));
    InMux I__10735 (
            .O(N__46568),
            .I(N__46560));
    LocalMux I__10734 (
            .O(N__46563),
            .I(N__46557));
    LocalMux I__10733 (
            .O(N__46560),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv12 I__10732 (
            .O(N__46557),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__10731 (
            .O(N__46552),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__10730 (
            .O(N__46549),
            .I(N__46542));
    InMux I__10729 (
            .O(N__46548),
            .I(N__46542));
    InMux I__10728 (
            .O(N__46547),
            .I(N__46539));
    LocalMux I__10727 (
            .O(N__46542),
            .I(N__46536));
    LocalMux I__10726 (
            .O(N__46539),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__10725 (
            .O(N__46536),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__10724 (
            .O(N__46531),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__10723 (
            .O(N__46528),
            .I(N__46525));
    InMux I__10722 (
            .O(N__46525),
            .I(N__46520));
    InMux I__10721 (
            .O(N__46524),
            .I(N__46517));
    InMux I__10720 (
            .O(N__46523),
            .I(N__46514));
    LocalMux I__10719 (
            .O(N__46520),
            .I(N__46511));
    LocalMux I__10718 (
            .O(N__46517),
            .I(N__46508));
    LocalMux I__10717 (
            .O(N__46514),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv12 I__10716 (
            .O(N__46511),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__10715 (
            .O(N__46508),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__10714 (
            .O(N__46501),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__10713 (
            .O(N__46498),
            .I(N__46493));
    InMux I__10712 (
            .O(N__46497),
            .I(N__46490));
    InMux I__10711 (
            .O(N__46496),
            .I(N__46487));
    LocalMux I__10710 (
            .O(N__46493),
            .I(N__46482));
    LocalMux I__10709 (
            .O(N__46490),
            .I(N__46482));
    LocalMux I__10708 (
            .O(N__46487),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__10707 (
            .O(N__46482),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__10706 (
            .O(N__46477),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__10705 (
            .O(N__46474),
            .I(N__46470));
    InMux I__10704 (
            .O(N__46473),
            .I(N__46467));
    LocalMux I__10703 (
            .O(N__46470),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__10702 (
            .O(N__46467),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__10701 (
            .O(N__46462),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__10700 (
            .O(N__46459),
            .I(N__46455));
    InMux I__10699 (
            .O(N__46458),
            .I(N__46452));
    LocalMux I__10698 (
            .O(N__46455),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__10697 (
            .O(N__46452),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__10696 (
            .O(N__46447),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__10695 (
            .O(N__46444),
            .I(N__46440));
    InMux I__10694 (
            .O(N__46443),
            .I(N__46437));
    LocalMux I__10693 (
            .O(N__46440),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__10692 (
            .O(N__46437),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__10691 (
            .O(N__46432),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__10690 (
            .O(N__46429),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__10689 (
            .O(N__46426),
            .I(bfn_18_12_0_));
    CascadeMux I__10688 (
            .O(N__46423),
            .I(N__46420));
    InMux I__10687 (
            .O(N__46420),
            .I(N__46415));
    InMux I__10686 (
            .O(N__46419),
            .I(N__46412));
    InMux I__10685 (
            .O(N__46418),
            .I(N__46409));
    LocalMux I__10684 (
            .O(N__46415),
            .I(N__46406));
    LocalMux I__10683 (
            .O(N__46412),
            .I(N__46403));
    LocalMux I__10682 (
            .O(N__46409),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__10681 (
            .O(N__46406),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv12 I__10680 (
            .O(N__46403),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__10679 (
            .O(N__46396),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__10678 (
            .O(N__46393),
            .I(N__46389));
    InMux I__10677 (
            .O(N__46392),
            .I(N__46385));
    InMux I__10676 (
            .O(N__46389),
            .I(N__46382));
    InMux I__10675 (
            .O(N__46388),
            .I(N__46379));
    LocalMux I__10674 (
            .O(N__46385),
            .I(N__46376));
    LocalMux I__10673 (
            .O(N__46382),
            .I(N__46373));
    LocalMux I__10672 (
            .O(N__46379),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__10671 (
            .O(N__46376),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv12 I__10670 (
            .O(N__46373),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__10669 (
            .O(N__46366),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    CascadeMux I__10668 (
            .O(N__46363),
            .I(N__46360));
    InMux I__10667 (
            .O(N__46360),
            .I(N__46355));
    InMux I__10666 (
            .O(N__46359),
            .I(N__46352));
    InMux I__10665 (
            .O(N__46358),
            .I(N__46349));
    LocalMux I__10664 (
            .O(N__46355),
            .I(N__46344));
    LocalMux I__10663 (
            .O(N__46352),
            .I(N__46344));
    LocalMux I__10662 (
            .O(N__46349),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__10661 (
            .O(N__46344),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__10660 (
            .O(N__46339),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__10659 (
            .O(N__46336),
            .I(N__46331));
    InMux I__10658 (
            .O(N__46335),
            .I(N__46328));
    InMux I__10657 (
            .O(N__46334),
            .I(N__46325));
    LocalMux I__10656 (
            .O(N__46331),
            .I(N__46320));
    LocalMux I__10655 (
            .O(N__46328),
            .I(N__46320));
    LocalMux I__10654 (
            .O(N__46325),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__10653 (
            .O(N__46320),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__10652 (
            .O(N__46315),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__10651 (
            .O(N__46312),
            .I(N__46308));
    InMux I__10650 (
            .O(N__46311),
            .I(N__46305));
    LocalMux I__10649 (
            .O(N__46308),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__10648 (
            .O(N__46305),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__10647 (
            .O(N__46300),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__10646 (
            .O(N__46297),
            .I(N__46293));
    InMux I__10645 (
            .O(N__46296),
            .I(N__46290));
    LocalMux I__10644 (
            .O(N__46293),
            .I(N__46287));
    LocalMux I__10643 (
            .O(N__46290),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__10642 (
            .O(N__46287),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__10641 (
            .O(N__46282),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__10640 (
            .O(N__46279),
            .I(N__46275));
    InMux I__10639 (
            .O(N__46278),
            .I(N__46272));
    LocalMux I__10638 (
            .O(N__46275),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__10637 (
            .O(N__46272),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__10636 (
            .O(N__46267),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__10635 (
            .O(N__46264),
            .I(N__46260));
    InMux I__10634 (
            .O(N__46263),
            .I(N__46257));
    LocalMux I__10633 (
            .O(N__46260),
            .I(N__46254));
    LocalMux I__10632 (
            .O(N__46257),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__10631 (
            .O(N__46254),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__10630 (
            .O(N__46249),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__10629 (
            .O(N__46246),
            .I(N__46242));
    InMux I__10628 (
            .O(N__46245),
            .I(N__46239));
    LocalMux I__10627 (
            .O(N__46242),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__10626 (
            .O(N__46239),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__10625 (
            .O(N__46234),
            .I(bfn_18_11_0_));
    InMux I__10624 (
            .O(N__46231),
            .I(N__46227));
    InMux I__10623 (
            .O(N__46230),
            .I(N__46224));
    LocalMux I__10622 (
            .O(N__46227),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__10621 (
            .O(N__46224),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__10620 (
            .O(N__46219),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__10619 (
            .O(N__46216),
            .I(N__46212));
    InMux I__10618 (
            .O(N__46215),
            .I(N__46209));
    LocalMux I__10617 (
            .O(N__46212),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__10616 (
            .O(N__46209),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10615 (
            .O(N__46204),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__10614 (
            .O(N__46201),
            .I(N__46197));
    InMux I__10613 (
            .O(N__46200),
            .I(N__46194));
    LocalMux I__10612 (
            .O(N__46197),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__10611 (
            .O(N__46194),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__10610 (
            .O(N__46189),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__10609 (
            .O(N__46186),
            .I(N__46182));
    InMux I__10608 (
            .O(N__46185),
            .I(N__46178));
    LocalMux I__10607 (
            .O(N__46182),
            .I(N__46175));
    InMux I__10606 (
            .O(N__46181),
            .I(N__46172));
    LocalMux I__10605 (
            .O(N__46178),
            .I(N__46169));
    Span4Mux_v I__10604 (
            .O(N__46175),
            .I(N__46163));
    LocalMux I__10603 (
            .O(N__46172),
            .I(N__46163));
    Span4Mux_v I__10602 (
            .O(N__46169),
            .I(N__46160));
    InMux I__10601 (
            .O(N__46168),
            .I(N__46157));
    Span4Mux_h I__10600 (
            .O(N__46163),
            .I(N__46154));
    Odrv4 I__10599 (
            .O(N__46160),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__10598 (
            .O(N__46157),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__10597 (
            .O(N__46154),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10596 (
            .O(N__46147),
            .I(N__46143));
    InMux I__10595 (
            .O(N__46146),
            .I(N__46140));
    LocalMux I__10594 (
            .O(N__46143),
            .I(N__46137));
    LocalMux I__10593 (
            .O(N__46140),
            .I(N__46133));
    Span4Mux_h I__10592 (
            .O(N__46137),
            .I(N__46130));
    InMux I__10591 (
            .O(N__46136),
            .I(N__46127));
    Span4Mux_h I__10590 (
            .O(N__46133),
            .I(N__46124));
    Span4Mux_v I__10589 (
            .O(N__46130),
            .I(N__46121));
    LocalMux I__10588 (
            .O(N__46127),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__10587 (
            .O(N__46124),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__10586 (
            .O(N__46121),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__10585 (
            .O(N__46114),
            .I(N__46111));
    LocalMux I__10584 (
            .O(N__46111),
            .I(N__46107));
    InMux I__10583 (
            .O(N__46110),
            .I(N__46104));
    Odrv4 I__10582 (
            .O(N__46107),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    LocalMux I__10581 (
            .O(N__46104),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    CascadeMux I__10580 (
            .O(N__46099),
            .I(N__46095));
    InMux I__10579 (
            .O(N__46098),
            .I(N__46092));
    InMux I__10578 (
            .O(N__46095),
            .I(N__46089));
    LocalMux I__10577 (
            .O(N__46092),
            .I(N__46086));
    LocalMux I__10576 (
            .O(N__46089),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    Odrv4 I__10575 (
            .O(N__46086),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__10574 (
            .O(N__46081),
            .I(N__46078));
    InMux I__10573 (
            .O(N__46078),
            .I(N__46075));
    LocalMux I__10572 (
            .O(N__46075),
            .I(N__46072));
    Span4Mux_v I__10571 (
            .O(N__46072),
            .I(N__46069));
    Odrv4 I__10570 (
            .O(N__46069),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__10569 (
            .O(N__46066),
            .I(N__46062));
    InMux I__10568 (
            .O(N__46065),
            .I(N__46059));
    LocalMux I__10567 (
            .O(N__46062),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    LocalMux I__10566 (
            .O(N__46059),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__10565 (
            .O(N__46054),
            .I(N__46050));
    InMux I__10564 (
            .O(N__46053),
            .I(N__46047));
    LocalMux I__10563 (
            .O(N__46050),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    LocalMux I__10562 (
            .O(N__46047),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__10561 (
            .O(N__46042),
            .I(N__46039));
    LocalMux I__10560 (
            .O(N__46039),
            .I(N__46036));
    Span4Mux_v I__10559 (
            .O(N__46036),
            .I(N__46033));
    Odrv4 I__10558 (
            .O(N__46033),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    CascadeMux I__10557 (
            .O(N__46030),
            .I(N__46026));
    InMux I__10556 (
            .O(N__46029),
            .I(N__46023));
    InMux I__10555 (
            .O(N__46026),
            .I(N__46020));
    LocalMux I__10554 (
            .O(N__46023),
            .I(N__46017));
    LocalMux I__10553 (
            .O(N__46020),
            .I(N__46011));
    Span4Mux_v I__10552 (
            .O(N__46017),
            .I(N__46011));
    InMux I__10551 (
            .O(N__46016),
            .I(N__46008));
    Odrv4 I__10550 (
            .O(N__46011),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__10549 (
            .O(N__46008),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__10548 (
            .O(N__46003),
            .I(N__45999));
    InMux I__10547 (
            .O(N__46002),
            .I(N__45996));
    LocalMux I__10546 (
            .O(N__45999),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__10545 (
            .O(N__45996),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__10544 (
            .O(N__45991),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__10543 (
            .O(N__45988),
            .I(N__45985));
    LocalMux I__10542 (
            .O(N__45985),
            .I(N__45982));
    Span4Mux_h I__10541 (
            .O(N__45982),
            .I(N__45979));
    Odrv4 I__10540 (
            .O(N__45979),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ));
    CascadeMux I__10539 (
            .O(N__45976),
            .I(N__45973));
    InMux I__10538 (
            .O(N__45973),
            .I(N__45969));
    InMux I__10537 (
            .O(N__45972),
            .I(N__45966));
    LocalMux I__10536 (
            .O(N__45969),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__10535 (
            .O(N__45966),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__10534 (
            .O(N__45961),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__10533 (
            .O(N__45958),
            .I(N__45954));
    InMux I__10532 (
            .O(N__45957),
            .I(N__45951));
    LocalMux I__10531 (
            .O(N__45954),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__10530 (
            .O(N__45951),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__10529 (
            .O(N__45946),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    CascadeMux I__10528 (
            .O(N__45943),
            .I(N__45938));
    InMux I__10527 (
            .O(N__45942),
            .I(N__45935));
    InMux I__10526 (
            .O(N__45941),
            .I(N__45932));
    InMux I__10525 (
            .O(N__45938),
            .I(N__45929));
    LocalMux I__10524 (
            .O(N__45935),
            .I(N__45925));
    LocalMux I__10523 (
            .O(N__45932),
            .I(N__45922));
    LocalMux I__10522 (
            .O(N__45929),
            .I(N__45919));
    InMux I__10521 (
            .O(N__45928),
            .I(N__45916));
    Span4Mux_h I__10520 (
            .O(N__45925),
            .I(N__45913));
    Span4Mux_v I__10519 (
            .O(N__45922),
            .I(N__45908));
    Span4Mux_v I__10518 (
            .O(N__45919),
            .I(N__45908));
    LocalMux I__10517 (
            .O(N__45916),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__10516 (
            .O(N__45913),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__10515 (
            .O(N__45908),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__10514 (
            .O(N__45901),
            .I(N__45897));
    InMux I__10513 (
            .O(N__45900),
            .I(N__45894));
    LocalMux I__10512 (
            .O(N__45897),
            .I(N__45890));
    LocalMux I__10511 (
            .O(N__45894),
            .I(N__45887));
    InMux I__10510 (
            .O(N__45893),
            .I(N__45884));
    Span4Mux_v I__10509 (
            .O(N__45890),
            .I(N__45881));
    Span4Mux_v I__10508 (
            .O(N__45887),
            .I(N__45878));
    LocalMux I__10507 (
            .O(N__45884),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__10506 (
            .O(N__45881),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__10505 (
            .O(N__45878),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__10504 (
            .O(N__45871),
            .I(N__45865));
    InMux I__10503 (
            .O(N__45870),
            .I(N__45865));
    LocalMux I__10502 (
            .O(N__45865),
            .I(N__45862));
    Odrv4 I__10501 (
            .O(N__45862),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__10500 (
            .O(N__45859),
            .I(N__45856));
    InMux I__10499 (
            .O(N__45856),
            .I(N__45850));
    InMux I__10498 (
            .O(N__45855),
            .I(N__45850));
    LocalMux I__10497 (
            .O(N__45850),
            .I(N__45847));
    Odrv4 I__10496 (
            .O(N__45847),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CEMux I__10495 (
            .O(N__45844),
            .I(N__45841));
    LocalMux I__10494 (
            .O(N__45841),
            .I(N__45837));
    CEMux I__10493 (
            .O(N__45840),
            .I(N__45829));
    Span4Mux_h I__10492 (
            .O(N__45837),
            .I(N__45820));
    CEMux I__10491 (
            .O(N__45836),
            .I(N__45817));
    CEMux I__10490 (
            .O(N__45835),
            .I(N__45811));
    InMux I__10489 (
            .O(N__45834),
            .I(N__45804));
    InMux I__10488 (
            .O(N__45833),
            .I(N__45804));
    InMux I__10487 (
            .O(N__45832),
            .I(N__45804));
    LocalMux I__10486 (
            .O(N__45829),
            .I(N__45801));
    InMux I__10485 (
            .O(N__45828),
            .I(N__45798));
    CEMux I__10484 (
            .O(N__45827),
            .I(N__45794));
    CEMux I__10483 (
            .O(N__45826),
            .I(N__45791));
    CEMux I__10482 (
            .O(N__45825),
            .I(N__45788));
    CEMux I__10481 (
            .O(N__45824),
            .I(N__45785));
    CEMux I__10480 (
            .O(N__45823),
            .I(N__45766));
    Span4Mux_v I__10479 (
            .O(N__45820),
            .I(N__45761));
    LocalMux I__10478 (
            .O(N__45817),
            .I(N__45761));
    InMux I__10477 (
            .O(N__45816),
            .I(N__45746));
    InMux I__10476 (
            .O(N__45815),
            .I(N__45746));
    InMux I__10475 (
            .O(N__45814),
            .I(N__45746));
    LocalMux I__10474 (
            .O(N__45811),
            .I(N__45743));
    LocalMux I__10473 (
            .O(N__45804),
            .I(N__45736));
    Span4Mux_h I__10472 (
            .O(N__45801),
            .I(N__45736));
    LocalMux I__10471 (
            .O(N__45798),
            .I(N__45736));
    CEMux I__10470 (
            .O(N__45797),
            .I(N__45733));
    LocalMux I__10469 (
            .O(N__45794),
            .I(N__45726));
    LocalMux I__10468 (
            .O(N__45791),
            .I(N__45726));
    LocalMux I__10467 (
            .O(N__45788),
            .I(N__45726));
    LocalMux I__10466 (
            .O(N__45785),
            .I(N__45723));
    InMux I__10465 (
            .O(N__45784),
            .I(N__45714));
    InMux I__10464 (
            .O(N__45783),
            .I(N__45714));
    InMux I__10463 (
            .O(N__45782),
            .I(N__45714));
    InMux I__10462 (
            .O(N__45781),
            .I(N__45714));
    InMux I__10461 (
            .O(N__45780),
            .I(N__45705));
    InMux I__10460 (
            .O(N__45779),
            .I(N__45705));
    InMux I__10459 (
            .O(N__45778),
            .I(N__45705));
    InMux I__10458 (
            .O(N__45777),
            .I(N__45705));
    InMux I__10457 (
            .O(N__45776),
            .I(N__45696));
    InMux I__10456 (
            .O(N__45775),
            .I(N__45696));
    InMux I__10455 (
            .O(N__45774),
            .I(N__45696));
    InMux I__10454 (
            .O(N__45773),
            .I(N__45696));
    InMux I__10453 (
            .O(N__45772),
            .I(N__45687));
    InMux I__10452 (
            .O(N__45771),
            .I(N__45687));
    InMux I__10451 (
            .O(N__45770),
            .I(N__45687));
    InMux I__10450 (
            .O(N__45769),
            .I(N__45687));
    LocalMux I__10449 (
            .O(N__45766),
            .I(N__45682));
    Span4Mux_h I__10448 (
            .O(N__45761),
            .I(N__45682));
    InMux I__10447 (
            .O(N__45760),
            .I(N__45673));
    InMux I__10446 (
            .O(N__45759),
            .I(N__45673));
    InMux I__10445 (
            .O(N__45758),
            .I(N__45673));
    InMux I__10444 (
            .O(N__45757),
            .I(N__45673));
    InMux I__10443 (
            .O(N__45756),
            .I(N__45664));
    InMux I__10442 (
            .O(N__45755),
            .I(N__45664));
    InMux I__10441 (
            .O(N__45754),
            .I(N__45664));
    InMux I__10440 (
            .O(N__45753),
            .I(N__45664));
    LocalMux I__10439 (
            .O(N__45746),
            .I(N__45657));
    Span4Mux_v I__10438 (
            .O(N__45743),
            .I(N__45657));
    Span4Mux_v I__10437 (
            .O(N__45736),
            .I(N__45657));
    LocalMux I__10436 (
            .O(N__45733),
            .I(N__45650));
    Sp12to4 I__10435 (
            .O(N__45726),
            .I(N__45650));
    Sp12to4 I__10434 (
            .O(N__45723),
            .I(N__45650));
    LocalMux I__10433 (
            .O(N__45714),
            .I(N__45639));
    LocalMux I__10432 (
            .O(N__45705),
            .I(N__45639));
    LocalMux I__10431 (
            .O(N__45696),
            .I(N__45639));
    LocalMux I__10430 (
            .O(N__45687),
            .I(N__45639));
    Span4Mux_v I__10429 (
            .O(N__45682),
            .I(N__45639));
    LocalMux I__10428 (
            .O(N__45673),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__10427 (
            .O(N__45664),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__10426 (
            .O(N__45657),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv12 I__10425 (
            .O(N__45650),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__10424 (
            .O(N__45639),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    CascadeMux I__10423 (
            .O(N__45628),
            .I(N__45625));
    InMux I__10422 (
            .O(N__45625),
            .I(N__45622));
    LocalMux I__10421 (
            .O(N__45622),
            .I(N__45619));
    Sp12to4 I__10420 (
            .O(N__45619),
            .I(N__45616));
    Odrv12 I__10419 (
            .O(N__45616),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    InMux I__10418 (
            .O(N__45613),
            .I(N__45610));
    LocalMux I__10417 (
            .O(N__45610),
            .I(N__45607));
    Span4Mux_h I__10416 (
            .O(N__45607),
            .I(N__45602));
    InMux I__10415 (
            .O(N__45606),
            .I(N__45599));
    InMux I__10414 (
            .O(N__45605),
            .I(N__45596));
    Span4Mux_v I__10413 (
            .O(N__45602),
            .I(N__45593));
    LocalMux I__10412 (
            .O(N__45599),
            .I(N__45590));
    LocalMux I__10411 (
            .O(N__45596),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv4 I__10410 (
            .O(N__45593),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv4 I__10409 (
            .O(N__45590),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__10408 (
            .O(N__45583),
            .I(N__45579));
    InMux I__10407 (
            .O(N__45582),
            .I(N__45575));
    LocalMux I__10406 (
            .O(N__45579),
            .I(N__45571));
    InMux I__10405 (
            .O(N__45578),
            .I(N__45568));
    LocalMux I__10404 (
            .O(N__45575),
            .I(N__45565));
    InMux I__10403 (
            .O(N__45574),
            .I(N__45562));
    Span4Mux_v I__10402 (
            .O(N__45571),
            .I(N__45557));
    LocalMux I__10401 (
            .O(N__45568),
            .I(N__45557));
    Span4Mux_h I__10400 (
            .O(N__45565),
            .I(N__45554));
    LocalMux I__10399 (
            .O(N__45562),
            .I(N__45551));
    Span4Mux_h I__10398 (
            .O(N__45557),
            .I(N__45548));
    Odrv4 I__10397 (
            .O(N__45554),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv12 I__10396 (
            .O(N__45551),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__10395 (
            .O(N__45548),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__10394 (
            .O(N__45541),
            .I(N__45538));
    LocalMux I__10393 (
            .O(N__45538),
            .I(N__45533));
    InMux I__10392 (
            .O(N__45537),
            .I(N__45530));
    InMux I__10391 (
            .O(N__45536),
            .I(N__45527));
    Span4Mux_h I__10390 (
            .O(N__45533),
            .I(N__45524));
    LocalMux I__10389 (
            .O(N__45530),
            .I(N__45521));
    LocalMux I__10388 (
            .O(N__45527),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__10387 (
            .O(N__45524),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__10386 (
            .O(N__45521),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__10385 (
            .O(N__45514),
            .I(N__45510));
    InMux I__10384 (
            .O(N__45513),
            .I(N__45506));
    LocalMux I__10383 (
            .O(N__45510),
            .I(N__45503));
    InMux I__10382 (
            .O(N__45509),
            .I(N__45499));
    LocalMux I__10381 (
            .O(N__45506),
            .I(N__45496));
    Span4Mux_v I__10380 (
            .O(N__45503),
            .I(N__45493));
    InMux I__10379 (
            .O(N__45502),
            .I(N__45490));
    LocalMux I__10378 (
            .O(N__45499),
            .I(N__45487));
    Span4Mux_v I__10377 (
            .O(N__45496),
            .I(N__45484));
    Odrv4 I__10376 (
            .O(N__45493),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__10375 (
            .O(N__45490),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__10374 (
            .O(N__45487),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__10373 (
            .O(N__45484),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__10372 (
            .O(N__45475),
            .I(N__45472));
    LocalMux I__10371 (
            .O(N__45472),
            .I(N__45468));
    InMux I__10370 (
            .O(N__45471),
            .I(N__45464));
    Span4Mux_v I__10369 (
            .O(N__45468),
            .I(N__45461));
    InMux I__10368 (
            .O(N__45467),
            .I(N__45458));
    LocalMux I__10367 (
            .O(N__45464),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__10366 (
            .O(N__45461),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__10365 (
            .O(N__45458),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__10364 (
            .O(N__45451),
            .I(N__45447));
    InMux I__10363 (
            .O(N__45450),
            .I(N__45443));
    LocalMux I__10362 (
            .O(N__45447),
            .I(N__45439));
    InMux I__10361 (
            .O(N__45446),
            .I(N__45436));
    LocalMux I__10360 (
            .O(N__45443),
            .I(N__45433));
    InMux I__10359 (
            .O(N__45442),
            .I(N__45430));
    Span4Mux_v I__10358 (
            .O(N__45439),
            .I(N__45427));
    LocalMux I__10357 (
            .O(N__45436),
            .I(N__45422));
    Span4Mux_v I__10356 (
            .O(N__45433),
            .I(N__45422));
    LocalMux I__10355 (
            .O(N__45430),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__10354 (
            .O(N__45427),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__10353 (
            .O(N__45422),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__10352 (
            .O(N__45415),
            .I(N__45412));
    InMux I__10351 (
            .O(N__45412),
            .I(N__45409));
    LocalMux I__10350 (
            .O(N__45409),
            .I(N__45406));
    Odrv4 I__10349 (
            .O(N__45406),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__10348 (
            .O(N__45403),
            .I(N__45400));
    LocalMux I__10347 (
            .O(N__45400),
            .I(N__45394));
    InMux I__10346 (
            .O(N__45399),
            .I(N__45391));
    InMux I__10345 (
            .O(N__45398),
            .I(N__45388));
    InMux I__10344 (
            .O(N__45397),
            .I(N__45385));
    Span4Mux_v I__10343 (
            .O(N__45394),
            .I(N__45378));
    LocalMux I__10342 (
            .O(N__45391),
            .I(N__45378));
    LocalMux I__10341 (
            .O(N__45388),
            .I(N__45378));
    LocalMux I__10340 (
            .O(N__45385),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__10339 (
            .O(N__45378),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__10338 (
            .O(N__45373),
            .I(N__45370));
    LocalMux I__10337 (
            .O(N__45370),
            .I(N__45366));
    InMux I__10336 (
            .O(N__45369),
            .I(N__45362));
    Span4Mux_v I__10335 (
            .O(N__45366),
            .I(N__45359));
    InMux I__10334 (
            .O(N__45365),
            .I(N__45356));
    LocalMux I__10333 (
            .O(N__45362),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__10332 (
            .O(N__45359),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__10331 (
            .O(N__45356),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__10330 (
            .O(N__45349),
            .I(N__45346));
    LocalMux I__10329 (
            .O(N__45346),
            .I(N__45343));
    Odrv4 I__10328 (
            .O(N__45343),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__10327 (
            .O(N__45340),
            .I(N__45337));
    LocalMux I__10326 (
            .O(N__45337),
            .I(N__45333));
    InMux I__10325 (
            .O(N__45336),
            .I(N__45329));
    Span4Mux_v I__10324 (
            .O(N__45333),
            .I(N__45326));
    InMux I__10323 (
            .O(N__45332),
            .I(N__45323));
    LocalMux I__10322 (
            .O(N__45329),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__10321 (
            .O(N__45326),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__10320 (
            .O(N__45323),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__10319 (
            .O(N__45316),
            .I(N__45313));
    LocalMux I__10318 (
            .O(N__45313),
            .I(N__45310));
    Odrv4 I__10317 (
            .O(N__45310),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__10316 (
            .O(N__45307),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__10315 (
            .O(N__45304),
            .I(N__45301));
    LocalMux I__10314 (
            .O(N__45301),
            .I(N__45297));
    InMux I__10313 (
            .O(N__45300),
            .I(N__45293));
    Span4Mux_v I__10312 (
            .O(N__45297),
            .I(N__45290));
    InMux I__10311 (
            .O(N__45296),
            .I(N__45287));
    LocalMux I__10310 (
            .O(N__45293),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__10309 (
            .O(N__45290),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__10308 (
            .O(N__45287),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__10307 (
            .O(N__45280),
            .I(N__45277));
    LocalMux I__10306 (
            .O(N__45277),
            .I(N__45274));
    Odrv4 I__10305 (
            .O(N__45274),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__10304 (
            .O(N__45271),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__10303 (
            .O(N__45268),
            .I(N__45264));
    InMux I__10302 (
            .O(N__45267),
            .I(N__45261));
    LocalMux I__10301 (
            .O(N__45264),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__10300 (
            .O(N__45261),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__10299 (
            .O(N__45256),
            .I(N__45253));
    LocalMux I__10298 (
            .O(N__45253),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__10297 (
            .O(N__45250),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__10296 (
            .O(N__45247),
            .I(N__45244));
    LocalMux I__10295 (
            .O(N__45244),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__10294 (
            .O(N__45241),
            .I(bfn_17_28_0_));
    InMux I__10293 (
            .O(N__45238),
            .I(N__45235));
    LocalMux I__10292 (
            .O(N__45235),
            .I(N__45231));
    InMux I__10291 (
            .O(N__45234),
            .I(N__45228));
    Span4Mux_s3_v I__10290 (
            .O(N__45231),
            .I(N__45225));
    LocalMux I__10289 (
            .O(N__45228),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__10288 (
            .O(N__45225),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__10287 (
            .O(N__45220),
            .I(N__45217));
    LocalMux I__10286 (
            .O(N__45217),
            .I(N__45214));
    Span4Mux_v I__10285 (
            .O(N__45214),
            .I(N__45211));
    Span4Mux_s2_v I__10284 (
            .O(N__45211),
            .I(N__45208));
    Odrv4 I__10283 (
            .O(N__45208),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__10282 (
            .O(N__45205),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__10281 (
            .O(N__45202),
            .I(N__45197));
    InMux I__10280 (
            .O(N__45201),
            .I(N__45194));
    InMux I__10279 (
            .O(N__45200),
            .I(N__45191));
    LocalMux I__10278 (
            .O(N__45197),
            .I(N__45188));
    LocalMux I__10277 (
            .O(N__45194),
            .I(N__45185));
    LocalMux I__10276 (
            .O(N__45191),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__10275 (
            .O(N__45188),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__10274 (
            .O(N__45185),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__10273 (
            .O(N__45178),
            .I(N__45175));
    LocalMux I__10272 (
            .O(N__45175),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__10271 (
            .O(N__45172),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__10270 (
            .O(N__45169),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__10269 (
            .O(N__45166),
            .I(N__45163));
    LocalMux I__10268 (
            .O(N__45163),
            .I(N__45160));
    Span4Mux_h I__10267 (
            .O(N__45160),
            .I(N__45157));
    Odrv4 I__10266 (
            .O(N__45157),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    CascadeMux I__10265 (
            .O(N__45154),
            .I(N__45150));
    InMux I__10264 (
            .O(N__45153),
            .I(N__45147));
    InMux I__10263 (
            .O(N__45150),
            .I(N__45144));
    LocalMux I__10262 (
            .O(N__45147),
            .I(N__45141));
    LocalMux I__10261 (
            .O(N__45144),
            .I(N__45138));
    Span4Mux_h I__10260 (
            .O(N__45141),
            .I(N__45135));
    Odrv4 I__10259 (
            .O(N__45138),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    Odrv4 I__10258 (
            .O(N__45135),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__10257 (
            .O(N__45130),
            .I(N__45125));
    InMux I__10256 (
            .O(N__45129),
            .I(N__45120));
    InMux I__10255 (
            .O(N__45128),
            .I(N__45120));
    LocalMux I__10254 (
            .O(N__45125),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__10253 (
            .O(N__45120),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__10252 (
            .O(N__45115),
            .I(N__45112));
    LocalMux I__10251 (
            .O(N__45112),
            .I(N__45109));
    Span4Mux_h I__10250 (
            .O(N__45109),
            .I(N__45106));
    Span4Mux_h I__10249 (
            .O(N__45106),
            .I(N__45103));
    Odrv4 I__10248 (
            .O(N__45103),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__10247 (
            .O(N__45100),
            .I(N__45097));
    LocalMux I__10246 (
            .O(N__45097),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__10245 (
            .O(N__45094),
            .I(N__45091));
    LocalMux I__10244 (
            .O(N__45091),
            .I(N__45088));
    Span4Mux_h I__10243 (
            .O(N__45088),
            .I(N__45085));
    Span4Mux_h I__10242 (
            .O(N__45085),
            .I(N__45082));
    Odrv4 I__10241 (
            .O(N__45082),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__10240 (
            .O(N__45079),
            .I(N__45076));
    LocalMux I__10239 (
            .O(N__45076),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__10238 (
            .O(N__45073),
            .I(N__45070));
    LocalMux I__10237 (
            .O(N__45070),
            .I(N__45067));
    Span4Mux_h I__10236 (
            .O(N__45067),
            .I(N__45064));
    Span4Mux_h I__10235 (
            .O(N__45064),
            .I(N__45061));
    Odrv4 I__10234 (
            .O(N__45061),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__10233 (
            .O(N__45058),
            .I(N__45055));
    LocalMux I__10232 (
            .O(N__45055),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__10231 (
            .O(N__45052),
            .I(N__45049));
    LocalMux I__10230 (
            .O(N__45049),
            .I(N__45046));
    Span4Mux_v I__10229 (
            .O(N__45046),
            .I(N__45043));
    Span4Mux_h I__10228 (
            .O(N__45043),
            .I(N__45040));
    Span4Mux_h I__10227 (
            .O(N__45040),
            .I(N__45037));
    Odrv4 I__10226 (
            .O(N__45037),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__10225 (
            .O(N__45034),
            .I(N__45031));
    LocalMux I__10224 (
            .O(N__45031),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__10223 (
            .O(N__45028),
            .I(N__45025));
    LocalMux I__10222 (
            .O(N__45025),
            .I(N__45022));
    Span4Mux_v I__10221 (
            .O(N__45022),
            .I(N__45019));
    Span4Mux_h I__10220 (
            .O(N__45019),
            .I(N__45016));
    Span4Mux_h I__10219 (
            .O(N__45016),
            .I(N__45013));
    Odrv4 I__10218 (
            .O(N__45013),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__10217 (
            .O(N__45010),
            .I(N__45007));
    LocalMux I__10216 (
            .O(N__45007),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__10215 (
            .O(N__45004),
            .I(N__45001));
    LocalMux I__10214 (
            .O(N__45001),
            .I(N__44998));
    Odrv12 I__10213 (
            .O(N__44998),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__10212 (
            .O(N__44995),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    CascadeMux I__10211 (
            .O(N__44992),
            .I(N__44986));
    CascadeMux I__10210 (
            .O(N__44991),
            .I(N__44980));
    CascadeMux I__10209 (
            .O(N__44990),
            .I(N__44977));
    CascadeMux I__10208 (
            .O(N__44989),
            .I(N__44973));
    InMux I__10207 (
            .O(N__44986),
            .I(N__44968));
    InMux I__10206 (
            .O(N__44985),
            .I(N__44961));
    InMux I__10205 (
            .O(N__44984),
            .I(N__44961));
    InMux I__10204 (
            .O(N__44983),
            .I(N__44961));
    InMux I__10203 (
            .O(N__44980),
            .I(N__44956));
    InMux I__10202 (
            .O(N__44977),
            .I(N__44956));
    InMux I__10201 (
            .O(N__44976),
            .I(N__44953));
    InMux I__10200 (
            .O(N__44973),
            .I(N__44950));
    CascadeMux I__10199 (
            .O(N__44972),
            .I(N__44946));
    InMux I__10198 (
            .O(N__44971),
            .I(N__44942));
    LocalMux I__10197 (
            .O(N__44968),
            .I(N__44937));
    LocalMux I__10196 (
            .O(N__44961),
            .I(N__44937));
    LocalMux I__10195 (
            .O(N__44956),
            .I(N__44934));
    LocalMux I__10194 (
            .O(N__44953),
            .I(N__44929));
    LocalMux I__10193 (
            .O(N__44950),
            .I(N__44929));
    InMux I__10192 (
            .O(N__44949),
            .I(N__44926));
    InMux I__10191 (
            .O(N__44946),
            .I(N__44921));
    InMux I__10190 (
            .O(N__44945),
            .I(N__44921));
    LocalMux I__10189 (
            .O(N__44942),
            .I(N__44918));
    Span4Mux_h I__10188 (
            .O(N__44937),
            .I(N__44913));
    Span4Mux_h I__10187 (
            .O(N__44934),
            .I(N__44913));
    Span4Mux_h I__10186 (
            .O(N__44929),
            .I(N__44908));
    LocalMux I__10185 (
            .O(N__44926),
            .I(N__44908));
    LocalMux I__10184 (
            .O(N__44921),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__10183 (
            .O(N__44918),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__10182 (
            .O(N__44913),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__10181 (
            .O(N__44908),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__10180 (
            .O(N__44899),
            .I(N__44895));
    InMux I__10179 (
            .O(N__44898),
            .I(N__44892));
    LocalMux I__10178 (
            .O(N__44895),
            .I(N__44889));
    LocalMux I__10177 (
            .O(N__44892),
            .I(N__44886));
    Span4Mux_v I__10176 (
            .O(N__44889),
            .I(N__44883));
    Span4Mux_h I__10175 (
            .O(N__44886),
            .I(N__44880));
    Span4Mux_h I__10174 (
            .O(N__44883),
            .I(N__44877));
    Span4Mux_h I__10173 (
            .O(N__44880),
            .I(N__44874));
    Span4Mux_h I__10172 (
            .O(N__44877),
            .I(N__44871));
    Odrv4 I__10171 (
            .O(N__44874),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__10170 (
            .O(N__44871),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__10169 (
            .O(N__44866),
            .I(N__44863));
    LocalMux I__10168 (
            .O(N__44863),
            .I(N__44860));
    Span4Mux_h I__10167 (
            .O(N__44860),
            .I(N__44857));
    Odrv4 I__10166 (
            .O(N__44857),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__10165 (
            .O(N__44854),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    CascadeMux I__10164 (
            .O(N__44851),
            .I(N__44848));
    InMux I__10163 (
            .O(N__44848),
            .I(N__44845));
    LocalMux I__10162 (
            .O(N__44845),
            .I(N__44841));
    InMux I__10161 (
            .O(N__44844),
            .I(N__44837));
    Span4Mux_h I__10160 (
            .O(N__44841),
            .I(N__44834));
    InMux I__10159 (
            .O(N__44840),
            .I(N__44831));
    LocalMux I__10158 (
            .O(N__44837),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__10157 (
            .O(N__44834),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__10156 (
            .O(N__44831),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__10155 (
            .O(N__44824),
            .I(N__44821));
    LocalMux I__10154 (
            .O(N__44821),
            .I(N__44818));
    Odrv12 I__10153 (
            .O(N__44818),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__10152 (
            .O(N__44815),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__10151 (
            .O(N__44812),
            .I(N__44808));
    InMux I__10150 (
            .O(N__44811),
            .I(N__44805));
    LocalMux I__10149 (
            .O(N__44808),
            .I(N__44799));
    LocalMux I__10148 (
            .O(N__44805),
            .I(N__44799));
    InMux I__10147 (
            .O(N__44804),
            .I(N__44796));
    Span4Mux_s3_v I__10146 (
            .O(N__44799),
            .I(N__44792));
    LocalMux I__10145 (
            .O(N__44796),
            .I(N__44789));
    InMux I__10144 (
            .O(N__44795),
            .I(N__44786));
    Span4Mux_h I__10143 (
            .O(N__44792),
            .I(N__44783));
    Span4Mux_v I__10142 (
            .O(N__44789),
            .I(N__44778));
    LocalMux I__10141 (
            .O(N__44786),
            .I(N__44778));
    Sp12to4 I__10140 (
            .O(N__44783),
            .I(N__44774));
    Span4Mux_v I__10139 (
            .O(N__44778),
            .I(N__44771));
    InMux I__10138 (
            .O(N__44777),
            .I(N__44768));
    Span12Mux_v I__10137 (
            .O(N__44774),
            .I(N__44765));
    Sp12to4 I__10136 (
            .O(N__44771),
            .I(N__44762));
    LocalMux I__10135 (
            .O(N__44768),
            .I(N__44759));
    Span12Mux_v I__10134 (
            .O(N__44765),
            .I(N__44756));
    Span12Mux_s7_h I__10133 (
            .O(N__44762),
            .I(N__44751));
    Sp12to4 I__10132 (
            .O(N__44759),
            .I(N__44751));
    Span12Mux_h I__10131 (
            .O(N__44756),
            .I(N__44748));
    Span12Mux_v I__10130 (
            .O(N__44751),
            .I(N__44745));
    Odrv12 I__10129 (
            .O(N__44748),
            .I(start_stop_c));
    Odrv12 I__10128 (
            .O(N__44745),
            .I(start_stop_c));
    CascadeMux I__10127 (
            .O(N__44740),
            .I(N__44736));
    InMux I__10126 (
            .O(N__44739),
            .I(N__44730));
    InMux I__10125 (
            .O(N__44736),
            .I(N__44725));
    InMux I__10124 (
            .O(N__44735),
            .I(N__44722));
    InMux I__10123 (
            .O(N__44734),
            .I(N__44717));
    InMux I__10122 (
            .O(N__44733),
            .I(N__44717));
    LocalMux I__10121 (
            .O(N__44730),
            .I(N__44714));
    InMux I__10120 (
            .O(N__44729),
            .I(N__44708));
    InMux I__10119 (
            .O(N__44728),
            .I(N__44708));
    LocalMux I__10118 (
            .O(N__44725),
            .I(N__44705));
    LocalMux I__10117 (
            .O(N__44722),
            .I(N__44700));
    LocalMux I__10116 (
            .O(N__44717),
            .I(N__44700));
    Span4Mux_h I__10115 (
            .O(N__44714),
            .I(N__44697));
    InMux I__10114 (
            .O(N__44713),
            .I(N__44694));
    LocalMux I__10113 (
            .O(N__44708),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__10112 (
            .O(N__44705),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__10111 (
            .O(N__44700),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__10110 (
            .O(N__44697),
            .I(phase_controller_inst1_state_4));
    LocalMux I__10109 (
            .O(N__44694),
            .I(phase_controller_inst1_state_4));
    InMux I__10108 (
            .O(N__44683),
            .I(N__44679));
    InMux I__10107 (
            .O(N__44682),
            .I(N__44676));
    LocalMux I__10106 (
            .O(N__44679),
            .I(state_ns_i_a3_1));
    LocalMux I__10105 (
            .O(N__44676),
            .I(state_ns_i_a3_1));
    InMux I__10104 (
            .O(N__44671),
            .I(N__44667));
    InMux I__10103 (
            .O(N__44670),
            .I(N__44664));
    LocalMux I__10102 (
            .O(N__44667),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__10101 (
            .O(N__44664),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__10100 (
            .O(N__44659),
            .I(N__44654));
    InMux I__10099 (
            .O(N__44658),
            .I(N__44651));
    InMux I__10098 (
            .O(N__44657),
            .I(N__44648));
    LocalMux I__10097 (
            .O(N__44654),
            .I(N__44643));
    LocalMux I__10096 (
            .O(N__44651),
            .I(N__44643));
    LocalMux I__10095 (
            .O(N__44648),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__10094 (
            .O(N__44643),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__10093 (
            .O(N__44638),
            .I(N__44632));
    InMux I__10092 (
            .O(N__44637),
            .I(N__44632));
    LocalMux I__10091 (
            .O(N__44632),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__10090 (
            .O(N__44629),
            .I(N__44626));
    LocalMux I__10089 (
            .O(N__44626),
            .I(N__44623));
    Span4Mux_v I__10088 (
            .O(N__44623),
            .I(N__44620));
    Span4Mux_h I__10087 (
            .O(N__44620),
            .I(N__44617));
    Span4Mux_h I__10086 (
            .O(N__44617),
            .I(N__44614));
    Odrv4 I__10085 (
            .O(N__44614),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__10084 (
            .O(N__44611),
            .I(N__44608));
    LocalMux I__10083 (
            .O(N__44608),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__10082 (
            .O(N__44605),
            .I(N__44602));
    LocalMux I__10081 (
            .O(N__44602),
            .I(N__44599));
    Span4Mux_v I__10080 (
            .O(N__44599),
            .I(N__44596));
    Span4Mux_h I__10079 (
            .O(N__44596),
            .I(N__44593));
    Span4Mux_h I__10078 (
            .O(N__44593),
            .I(N__44590));
    Odrv4 I__10077 (
            .O(N__44590),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__10076 (
            .O(N__44587),
            .I(N__44584));
    LocalMux I__10075 (
            .O(N__44584),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__10074 (
            .O(N__44581),
            .I(N__44578));
    LocalMux I__10073 (
            .O(N__44578),
            .I(N__44575));
    Span4Mux_h I__10072 (
            .O(N__44575),
            .I(N__44572));
    Span4Mux_h I__10071 (
            .O(N__44572),
            .I(N__44569));
    Odrv4 I__10070 (
            .O(N__44569),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__10069 (
            .O(N__44566),
            .I(N__44563));
    LocalMux I__10068 (
            .O(N__44563),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__10067 (
            .O(N__44560),
            .I(N__44557));
    LocalMux I__10066 (
            .O(N__44557),
            .I(N__44554));
    Span12Mux_h I__10065 (
            .O(N__44554),
            .I(N__44551));
    Odrv12 I__10064 (
            .O(N__44551),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__10063 (
            .O(N__44548),
            .I(N__44545));
    LocalMux I__10062 (
            .O(N__44545),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__10061 (
            .O(N__44542),
            .I(N__44539));
    LocalMux I__10060 (
            .O(N__44539),
            .I(N__44536));
    Span12Mux_s7_v I__10059 (
            .O(N__44536),
            .I(N__44533));
    Odrv12 I__10058 (
            .O(N__44533),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__10057 (
            .O(N__44530),
            .I(N__44527));
    LocalMux I__10056 (
            .O(N__44527),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__10055 (
            .O(N__44524),
            .I(N__44521));
    LocalMux I__10054 (
            .O(N__44521),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    CascadeMux I__10053 (
            .O(N__44518),
            .I(N__44515));
    InMux I__10052 (
            .O(N__44515),
            .I(N__44512));
    LocalMux I__10051 (
            .O(N__44512),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    InMux I__10050 (
            .O(N__44509),
            .I(N__44506));
    LocalMux I__10049 (
            .O(N__44506),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    CascadeMux I__10048 (
            .O(N__44503),
            .I(N__44500));
    InMux I__10047 (
            .O(N__44500),
            .I(N__44497));
    LocalMux I__10046 (
            .O(N__44497),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    InMux I__10045 (
            .O(N__44494),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__10044 (
            .O(N__44491),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    IoInMux I__10043 (
            .O(N__44488),
            .I(N__44485));
    LocalMux I__10042 (
            .O(N__44485),
            .I(N__44482));
    Span4Mux_s3_v I__10041 (
            .O(N__44482),
            .I(N__44479));
    Span4Mux_v I__10040 (
            .O(N__44479),
            .I(N__44476));
    Span4Mux_v I__10039 (
            .O(N__44476),
            .I(N__44472));
    InMux I__10038 (
            .O(N__44475),
            .I(N__44469));
    Odrv4 I__10037 (
            .O(N__44472),
            .I(test_c));
    LocalMux I__10036 (
            .O(N__44469),
            .I(test_c));
    CascadeMux I__10035 (
            .O(N__44464),
            .I(N__44461));
    InMux I__10034 (
            .O(N__44461),
            .I(N__44458));
    LocalMux I__10033 (
            .O(N__44458),
            .I(N__44455));
    Odrv12 I__10032 (
            .O(N__44455),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__10031 (
            .O(N__44452),
            .I(N__44449));
    LocalMux I__10030 (
            .O(N__44449),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__10029 (
            .O(N__44446),
            .I(N__44443));
    InMux I__10028 (
            .O(N__44443),
            .I(N__44440));
    LocalMux I__10027 (
            .O(N__44440),
            .I(N__44437));
    Odrv12 I__10026 (
            .O(N__44437),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__10025 (
            .O(N__44434),
            .I(N__44431));
    LocalMux I__10024 (
            .O(N__44431),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__10023 (
            .O(N__44428),
            .I(N__44425));
    InMux I__10022 (
            .O(N__44425),
            .I(N__44422));
    LocalMux I__10021 (
            .O(N__44422),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__10020 (
            .O(N__44419),
            .I(N__44416));
    LocalMux I__10019 (
            .O(N__44416),
            .I(N__44413));
    Odrv12 I__10018 (
            .O(N__44413),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__10017 (
            .O(N__44410),
            .I(N__44407));
    InMux I__10016 (
            .O(N__44407),
            .I(N__44404));
    LocalMux I__10015 (
            .O(N__44404),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__10014 (
            .O(N__44401),
            .I(N__44398));
    LocalMux I__10013 (
            .O(N__44398),
            .I(N__44395));
    Odrv12 I__10012 (
            .O(N__44395),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__10011 (
            .O(N__44392),
            .I(N__44389));
    LocalMux I__10010 (
            .O(N__44389),
            .I(N__44386));
    Odrv12 I__10009 (
            .O(N__44386),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    CascadeMux I__10008 (
            .O(N__44383),
            .I(N__44380));
    InMux I__10007 (
            .O(N__44380),
            .I(N__44377));
    LocalMux I__10006 (
            .O(N__44377),
            .I(N__44374));
    Odrv12 I__10005 (
            .O(N__44374),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__10004 (
            .O(N__44371),
            .I(N__44368));
    LocalMux I__10003 (
            .O(N__44368),
            .I(N__44365));
    Span4Mux_v I__10002 (
            .O(N__44365),
            .I(N__44362));
    Odrv4 I__10001 (
            .O(N__44362),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__10000 (
            .O(N__44359),
            .I(N__44356));
    InMux I__9999 (
            .O(N__44356),
            .I(N__44353));
    LocalMux I__9998 (
            .O(N__44353),
            .I(N__44350));
    Odrv4 I__9997 (
            .O(N__44350),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__9996 (
            .O(N__44347),
            .I(N__44344));
    InMux I__9995 (
            .O(N__44344),
            .I(N__44341));
    LocalMux I__9994 (
            .O(N__44341),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__9993 (
            .O(N__44338),
            .I(N__44335));
    LocalMux I__9992 (
            .O(N__44335),
            .I(N__44332));
    Odrv4 I__9991 (
            .O(N__44332),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__9990 (
            .O(N__44329),
            .I(N__44326));
    InMux I__9989 (
            .O(N__44326),
            .I(N__44323));
    LocalMux I__9988 (
            .O(N__44323),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__9987 (
            .O(N__44320),
            .I(N__44317));
    LocalMux I__9986 (
            .O(N__44317),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__9985 (
            .O(N__44314),
            .I(N__44311));
    InMux I__9984 (
            .O(N__44311),
            .I(N__44308));
    LocalMux I__9983 (
            .O(N__44308),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__9982 (
            .O(N__44305),
            .I(N__44302));
    LocalMux I__9981 (
            .O(N__44302),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__9980 (
            .O(N__44299),
            .I(N__44296));
    InMux I__9979 (
            .O(N__44296),
            .I(N__44293));
    LocalMux I__9978 (
            .O(N__44293),
            .I(N__44290));
    Odrv4 I__9977 (
            .O(N__44290),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__9976 (
            .O(N__44287),
            .I(N__44284));
    LocalMux I__9975 (
            .O(N__44284),
            .I(N__44281));
    Odrv12 I__9974 (
            .O(N__44281),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__9973 (
            .O(N__44278),
            .I(N__44275));
    InMux I__9972 (
            .O(N__44275),
            .I(N__44272));
    LocalMux I__9971 (
            .O(N__44272),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__9970 (
            .O(N__44269),
            .I(N__44266));
    LocalMux I__9969 (
            .O(N__44266),
            .I(N__44263));
    Odrv4 I__9968 (
            .O(N__44263),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__9967 (
            .O(N__44260),
            .I(N__44257));
    InMux I__9966 (
            .O(N__44257),
            .I(N__44254));
    LocalMux I__9965 (
            .O(N__44254),
            .I(N__44251));
    Odrv4 I__9964 (
            .O(N__44251),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__9963 (
            .O(N__44248),
            .I(N__44245));
    LocalMux I__9962 (
            .O(N__44245),
            .I(N__44242));
    Span4Mux_v I__9961 (
            .O(N__44242),
            .I(N__44239));
    Odrv4 I__9960 (
            .O(N__44239),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__9959 (
            .O(N__44236),
            .I(N__44233));
    InMux I__9958 (
            .O(N__44233),
            .I(N__44230));
    LocalMux I__9957 (
            .O(N__44230),
            .I(N__44227));
    Odrv4 I__9956 (
            .O(N__44227),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__9955 (
            .O(N__44224),
            .I(N__44220));
    InMux I__9954 (
            .O(N__44223),
            .I(N__44217));
    LocalMux I__9953 (
            .O(N__44220),
            .I(N__44212));
    LocalMux I__9952 (
            .O(N__44217),
            .I(N__44209));
    InMux I__9951 (
            .O(N__44216),
            .I(N__44204));
    InMux I__9950 (
            .O(N__44215),
            .I(N__44204));
    Span4Mux_h I__9949 (
            .O(N__44212),
            .I(N__44201));
    Span4Mux_h I__9948 (
            .O(N__44209),
            .I(N__44198));
    LocalMux I__9947 (
            .O(N__44204),
            .I(N__44195));
    Odrv4 I__9946 (
            .O(N__44201),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv4 I__9945 (
            .O(N__44198),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv12 I__9944 (
            .O(N__44195),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__9943 (
            .O(N__44188),
            .I(N__44183));
    InMux I__9942 (
            .O(N__44187),
            .I(N__44180));
    InMux I__9941 (
            .O(N__44186),
            .I(N__44177));
    LocalMux I__9940 (
            .O(N__44183),
            .I(N__44172));
    LocalMux I__9939 (
            .O(N__44180),
            .I(N__44172));
    LocalMux I__9938 (
            .O(N__44177),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    Odrv4 I__9937 (
            .O(N__44172),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__9936 (
            .O(N__44167),
            .I(N__44164));
    LocalMux I__9935 (
            .O(N__44164),
            .I(N__44160));
    InMux I__9934 (
            .O(N__44163),
            .I(N__44156));
    Span4Mux_v I__9933 (
            .O(N__44160),
            .I(N__44153));
    InMux I__9932 (
            .O(N__44159),
            .I(N__44150));
    LocalMux I__9931 (
            .O(N__44156),
            .I(N__44147));
    Span4Mux_h I__9930 (
            .O(N__44153),
            .I(N__44144));
    LocalMux I__9929 (
            .O(N__44150),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    Odrv12 I__9928 (
            .O(N__44147),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    Odrv4 I__9927 (
            .O(N__44144),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    CascadeMux I__9926 (
            .O(N__44137),
            .I(N__44132));
    InMux I__9925 (
            .O(N__44136),
            .I(N__44128));
    InMux I__9924 (
            .O(N__44135),
            .I(N__44125));
    InMux I__9923 (
            .O(N__44132),
            .I(N__44122));
    InMux I__9922 (
            .O(N__44131),
            .I(N__44119));
    LocalMux I__9921 (
            .O(N__44128),
            .I(N__44116));
    LocalMux I__9920 (
            .O(N__44125),
            .I(N__44113));
    LocalMux I__9919 (
            .O(N__44122),
            .I(N__44110));
    LocalMux I__9918 (
            .O(N__44119),
            .I(N__44101));
    Span4Mux_v I__9917 (
            .O(N__44116),
            .I(N__44101));
    Span4Mux_v I__9916 (
            .O(N__44113),
            .I(N__44101));
    Span4Mux_v I__9915 (
            .O(N__44110),
            .I(N__44101));
    Odrv4 I__9914 (
            .O(N__44101),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__9913 (
            .O(N__44098),
            .I(N__44095));
    LocalMux I__9912 (
            .O(N__44095),
            .I(N__44092));
    Span4Mux_h I__9911 (
            .O(N__44092),
            .I(N__44088));
    InMux I__9910 (
            .O(N__44091),
            .I(N__44084));
    Span4Mux_v I__9909 (
            .O(N__44088),
            .I(N__44081));
    InMux I__9908 (
            .O(N__44087),
            .I(N__44078));
    LocalMux I__9907 (
            .O(N__44084),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__9906 (
            .O(N__44081),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__9905 (
            .O(N__44078),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__9904 (
            .O(N__44071),
            .I(N__44066));
    InMux I__9903 (
            .O(N__44070),
            .I(N__44062));
    InMux I__9902 (
            .O(N__44069),
            .I(N__44059));
    LocalMux I__9901 (
            .O(N__44066),
            .I(N__44056));
    InMux I__9900 (
            .O(N__44065),
            .I(N__44053));
    LocalMux I__9899 (
            .O(N__44062),
            .I(N__44050));
    LocalMux I__9898 (
            .O(N__44059),
            .I(N__44047));
    Span4Mux_v I__9897 (
            .O(N__44056),
            .I(N__44042));
    LocalMux I__9896 (
            .O(N__44053),
            .I(N__44042));
    Odrv4 I__9895 (
            .O(N__44050),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__9894 (
            .O(N__44047),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__9893 (
            .O(N__44042),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__9892 (
            .O(N__44035),
            .I(N__44031));
    InMux I__9891 (
            .O(N__44034),
            .I(N__44028));
    LocalMux I__9890 (
            .O(N__44031),
            .I(N__44025));
    LocalMux I__9889 (
            .O(N__44028),
            .I(N__44021));
    Span4Mux_h I__9888 (
            .O(N__44025),
            .I(N__44018));
    InMux I__9887 (
            .O(N__44024),
            .I(N__44015));
    Span12Mux_h I__9886 (
            .O(N__44021),
            .I(N__44012));
    Span4Mux_v I__9885 (
            .O(N__44018),
            .I(N__44009));
    LocalMux I__9884 (
            .O(N__44015),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv12 I__9883 (
            .O(N__44012),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__9882 (
            .O(N__44009),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__9881 (
            .O(N__44002),
            .I(N__43997));
    InMux I__9880 (
            .O(N__44001),
            .I(N__43994));
    InMux I__9879 (
            .O(N__44000),
            .I(N__43991));
    LocalMux I__9878 (
            .O(N__43997),
            .I(N__43987));
    LocalMux I__9877 (
            .O(N__43994),
            .I(N__43984));
    LocalMux I__9876 (
            .O(N__43991),
            .I(N__43981));
    InMux I__9875 (
            .O(N__43990),
            .I(N__43978));
    Span4Mux_h I__9874 (
            .O(N__43987),
            .I(N__43973));
    Span4Mux_v I__9873 (
            .O(N__43984),
            .I(N__43973));
    Span4Mux_v I__9872 (
            .O(N__43981),
            .I(N__43970));
    LocalMux I__9871 (
            .O(N__43978),
            .I(N__43967));
    Odrv4 I__9870 (
            .O(N__43973),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__9869 (
            .O(N__43970),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__9868 (
            .O(N__43967),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    CascadeMux I__9867 (
            .O(N__43960),
            .I(N__43957));
    InMux I__9866 (
            .O(N__43957),
            .I(N__43954));
    LocalMux I__9865 (
            .O(N__43954),
            .I(N__43951));
    Span4Mux_v I__9864 (
            .O(N__43951),
            .I(N__43948));
    Odrv4 I__9863 (
            .O(N__43948),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    InMux I__9862 (
            .O(N__43945),
            .I(N__43942));
    LocalMux I__9861 (
            .O(N__43942),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__9860 (
            .O(N__43939),
            .I(N__43936));
    InMux I__9859 (
            .O(N__43936),
            .I(N__43933));
    LocalMux I__9858 (
            .O(N__43933),
            .I(N__43930));
    Odrv4 I__9857 (
            .O(N__43930),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__9856 (
            .O(N__43927),
            .I(N__43924));
    LocalMux I__9855 (
            .O(N__43924),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__9854 (
            .O(N__43921),
            .I(N__43918));
    LocalMux I__9853 (
            .O(N__43918),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__9852 (
            .O(N__43915),
            .I(N__43910));
    InMux I__9851 (
            .O(N__43914),
            .I(N__43907));
    InMux I__9850 (
            .O(N__43913),
            .I(N__43904));
    LocalMux I__9849 (
            .O(N__43910),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    LocalMux I__9848 (
            .O(N__43907),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    LocalMux I__9847 (
            .O(N__43904),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    CascadeMux I__9846 (
            .O(N__43897),
            .I(N__43892));
    CascadeMux I__9845 (
            .O(N__43896),
            .I(N__43889));
    CascadeMux I__9844 (
            .O(N__43895),
            .I(N__43885));
    InMux I__9843 (
            .O(N__43892),
            .I(N__43882));
    InMux I__9842 (
            .O(N__43889),
            .I(N__43879));
    InMux I__9841 (
            .O(N__43888),
            .I(N__43876));
    InMux I__9840 (
            .O(N__43885),
            .I(N__43873));
    LocalMux I__9839 (
            .O(N__43882),
            .I(N__43864));
    LocalMux I__9838 (
            .O(N__43879),
            .I(N__43864));
    LocalMux I__9837 (
            .O(N__43876),
            .I(N__43864));
    LocalMux I__9836 (
            .O(N__43873),
            .I(N__43864));
    Span4Mux_v I__9835 (
            .O(N__43864),
            .I(N__43861));
    Odrv4 I__9834 (
            .O(N__43861),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9833 (
            .O(N__43858),
            .I(N__43854));
    InMux I__9832 (
            .O(N__43857),
            .I(N__43850));
    LocalMux I__9831 (
            .O(N__43854),
            .I(N__43847));
    InMux I__9830 (
            .O(N__43853),
            .I(N__43843));
    LocalMux I__9829 (
            .O(N__43850),
            .I(N__43840));
    Span4Mux_h I__9828 (
            .O(N__43847),
            .I(N__43837));
    InMux I__9827 (
            .O(N__43846),
            .I(N__43834));
    LocalMux I__9826 (
            .O(N__43843),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__9825 (
            .O(N__43840),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__9824 (
            .O(N__43837),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__9823 (
            .O(N__43834),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__9822 (
            .O(N__43825),
            .I(N__43822));
    LocalMux I__9821 (
            .O(N__43822),
            .I(N__43818));
    InMux I__9820 (
            .O(N__43821),
            .I(N__43814));
    Span4Mux_h I__9819 (
            .O(N__43818),
            .I(N__43811));
    InMux I__9818 (
            .O(N__43817),
            .I(N__43808));
    LocalMux I__9817 (
            .O(N__43814),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv4 I__9816 (
            .O(N__43811),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    LocalMux I__9815 (
            .O(N__43808),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__9814 (
            .O(N__43801),
            .I(N__43796));
    InMux I__9813 (
            .O(N__43800),
            .I(N__43793));
    InMux I__9812 (
            .O(N__43799),
            .I(N__43790));
    LocalMux I__9811 (
            .O(N__43796),
            .I(N__43785));
    LocalMux I__9810 (
            .O(N__43793),
            .I(N__43785));
    LocalMux I__9809 (
            .O(N__43790),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv12 I__9808 (
            .O(N__43785),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__9807 (
            .O(N__43780),
            .I(N__43776));
    InMux I__9806 (
            .O(N__43779),
            .I(N__43773));
    LocalMux I__9805 (
            .O(N__43776),
            .I(N__43768));
    LocalMux I__9804 (
            .O(N__43773),
            .I(N__43765));
    InMux I__9803 (
            .O(N__43772),
            .I(N__43762));
    InMux I__9802 (
            .O(N__43771),
            .I(N__43759));
    Span4Mux_h I__9801 (
            .O(N__43768),
            .I(N__43754));
    Span4Mux_h I__9800 (
            .O(N__43765),
            .I(N__43754));
    LocalMux I__9799 (
            .O(N__43762),
            .I(N__43751));
    LocalMux I__9798 (
            .O(N__43759),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__9797 (
            .O(N__43754),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv12 I__9796 (
            .O(N__43751),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__9795 (
            .O(N__43744),
            .I(N__43740));
    InMux I__9794 (
            .O(N__43743),
            .I(N__43736));
    LocalMux I__9793 (
            .O(N__43740),
            .I(N__43733));
    InMux I__9792 (
            .O(N__43739),
            .I(N__43730));
    LocalMux I__9791 (
            .O(N__43736),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__9790 (
            .O(N__43733),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__9789 (
            .O(N__43730),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__9788 (
            .O(N__43723),
            .I(N__43718));
    InMux I__9787 (
            .O(N__43722),
            .I(N__43715));
    InMux I__9786 (
            .O(N__43721),
            .I(N__43712));
    LocalMux I__9785 (
            .O(N__43718),
            .I(N__43707));
    LocalMux I__9784 (
            .O(N__43715),
            .I(N__43707));
    LocalMux I__9783 (
            .O(N__43712),
            .I(N__43703));
    Span4Mux_v I__9782 (
            .O(N__43707),
            .I(N__43700));
    InMux I__9781 (
            .O(N__43706),
            .I(N__43697));
    Odrv4 I__9780 (
            .O(N__43703),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__9779 (
            .O(N__43700),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__9778 (
            .O(N__43697),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__9777 (
            .O(N__43690),
            .I(N__43686));
    InMux I__9776 (
            .O(N__43689),
            .I(N__43682));
    LocalMux I__9775 (
            .O(N__43686),
            .I(N__43679));
    InMux I__9774 (
            .O(N__43685),
            .I(N__43676));
    LocalMux I__9773 (
            .O(N__43682),
            .I(N__43671));
    Span4Mux_h I__9772 (
            .O(N__43679),
            .I(N__43671));
    LocalMux I__9771 (
            .O(N__43676),
            .I(N__43668));
    Odrv4 I__9770 (
            .O(N__43671),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    Odrv4 I__9769 (
            .O(N__43668),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__9768 (
            .O(N__43663),
            .I(N__43657));
    InMux I__9767 (
            .O(N__43662),
            .I(N__43654));
    InMux I__9766 (
            .O(N__43661),
            .I(N__43651));
    InMux I__9765 (
            .O(N__43660),
            .I(N__43648));
    LocalMux I__9764 (
            .O(N__43657),
            .I(N__43643));
    LocalMux I__9763 (
            .O(N__43654),
            .I(N__43643));
    LocalMux I__9762 (
            .O(N__43651),
            .I(N__43638));
    LocalMux I__9761 (
            .O(N__43648),
            .I(N__43638));
    Span4Mux_v I__9760 (
            .O(N__43643),
            .I(N__43635));
    Span4Mux_v I__9759 (
            .O(N__43638),
            .I(N__43632));
    Odrv4 I__9758 (
            .O(N__43635),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__9757 (
            .O(N__43632),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9756 (
            .O(N__43627),
            .I(N__43621));
    InMux I__9755 (
            .O(N__43626),
            .I(N__43621));
    LocalMux I__9754 (
            .O(N__43621),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__9753 (
            .O(N__43618),
            .I(N__43615));
    InMux I__9752 (
            .O(N__43615),
            .I(N__43609));
    InMux I__9751 (
            .O(N__43614),
            .I(N__43609));
    LocalMux I__9750 (
            .O(N__43609),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    InMux I__9749 (
            .O(N__43606),
            .I(N__43602));
    InMux I__9748 (
            .O(N__43605),
            .I(N__43599));
    LocalMux I__9747 (
            .O(N__43602),
            .I(N__43592));
    LocalMux I__9746 (
            .O(N__43599),
            .I(N__43592));
    InMux I__9745 (
            .O(N__43598),
            .I(N__43589));
    InMux I__9744 (
            .O(N__43597),
            .I(N__43586));
    Span4Mux_h I__9743 (
            .O(N__43592),
            .I(N__43583));
    LocalMux I__9742 (
            .O(N__43589),
            .I(N__43580));
    LocalMux I__9741 (
            .O(N__43586),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__9740 (
            .O(N__43583),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv12 I__9739 (
            .O(N__43580),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__9738 (
            .O(N__43573),
            .I(N__43569));
    InMux I__9737 (
            .O(N__43572),
            .I(N__43566));
    LocalMux I__9736 (
            .O(N__43569),
            .I(N__43559));
    LocalMux I__9735 (
            .O(N__43566),
            .I(N__43559));
    InMux I__9734 (
            .O(N__43565),
            .I(N__43556));
    InMux I__9733 (
            .O(N__43564),
            .I(N__43553));
    Span4Mux_v I__9732 (
            .O(N__43559),
            .I(N__43550));
    LocalMux I__9731 (
            .O(N__43556),
            .I(N__43547));
    LocalMux I__9730 (
            .O(N__43553),
            .I(N__43544));
    Span4Mux_h I__9729 (
            .O(N__43550),
            .I(N__43539));
    Span4Mux_v I__9728 (
            .O(N__43547),
            .I(N__43539));
    Odrv4 I__9727 (
            .O(N__43544),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__9726 (
            .O(N__43539),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__9725 (
            .O(N__43534),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ));
    InMux I__9724 (
            .O(N__43531),
            .I(N__43528));
    LocalMux I__9723 (
            .O(N__43528),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__9722 (
            .O(N__43525),
            .I(N__43522));
    LocalMux I__9721 (
            .O(N__43522),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__9720 (
            .O(N__43519),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    InMux I__9719 (
            .O(N__43516),
            .I(N__43513));
    LocalMux I__9718 (
            .O(N__43513),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    CascadeMux I__9717 (
            .O(N__43510),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__9716 (
            .O(N__43507),
            .I(N__43502));
    InMux I__9715 (
            .O(N__43506),
            .I(N__43499));
    InMux I__9714 (
            .O(N__43505),
            .I(N__43496));
    LocalMux I__9713 (
            .O(N__43502),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__9712 (
            .O(N__43499),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__9711 (
            .O(N__43496),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__9710 (
            .O(N__43489),
            .I(N__43485));
    InMux I__9709 (
            .O(N__43488),
            .I(N__43482));
    LocalMux I__9708 (
            .O(N__43485),
            .I(N__43476));
    LocalMux I__9707 (
            .O(N__43482),
            .I(N__43476));
    InMux I__9706 (
            .O(N__43481),
            .I(N__43473));
    Span4Mux_v I__9705 (
            .O(N__43476),
            .I(N__43467));
    LocalMux I__9704 (
            .O(N__43473),
            .I(N__43467));
    InMux I__9703 (
            .O(N__43472),
            .I(N__43464));
    Span4Mux_h I__9702 (
            .O(N__43467),
            .I(N__43461));
    LocalMux I__9701 (
            .O(N__43464),
            .I(N__43458));
    Odrv4 I__9700 (
            .O(N__43461),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv12 I__9699 (
            .O(N__43458),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__9698 (
            .O(N__43453),
            .I(N__43450));
    LocalMux I__9697 (
            .O(N__43450),
            .I(N__43445));
    InMux I__9696 (
            .O(N__43449),
            .I(N__43442));
    InMux I__9695 (
            .O(N__43448),
            .I(N__43439));
    Span4Mux_h I__9694 (
            .O(N__43445),
            .I(N__43436));
    LocalMux I__9693 (
            .O(N__43442),
            .I(N__43433));
    LocalMux I__9692 (
            .O(N__43439),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__9691 (
            .O(N__43436),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv12 I__9690 (
            .O(N__43433),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__9689 (
            .O(N__43426),
            .I(N__43423));
    LocalMux I__9688 (
            .O(N__43423),
            .I(N__43419));
    InMux I__9687 (
            .O(N__43422),
            .I(N__43416));
    Span4Mux_v I__9686 (
            .O(N__43419),
            .I(N__43409));
    LocalMux I__9685 (
            .O(N__43416),
            .I(N__43409));
    InMux I__9684 (
            .O(N__43415),
            .I(N__43406));
    InMux I__9683 (
            .O(N__43414),
            .I(N__43403));
    Span4Mux_h I__9682 (
            .O(N__43409),
            .I(N__43398));
    LocalMux I__9681 (
            .O(N__43406),
            .I(N__43398));
    LocalMux I__9680 (
            .O(N__43403),
            .I(N__43395));
    Odrv4 I__9679 (
            .O(N__43398),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv12 I__9678 (
            .O(N__43395),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    CascadeMux I__9677 (
            .O(N__43390),
            .I(N__43387));
    InMux I__9676 (
            .O(N__43387),
            .I(N__43384));
    LocalMux I__9675 (
            .O(N__43384),
            .I(N__43381));
    Span4Mux_v I__9674 (
            .O(N__43381),
            .I(N__43378));
    Sp12to4 I__9673 (
            .O(N__43378),
            .I(N__43375));
    Span12Mux_h I__9672 (
            .O(N__43375),
            .I(N__43372));
    Odrv12 I__9671 (
            .O(N__43372),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__9670 (
            .O(N__43369),
            .I(N__43366));
    LocalMux I__9669 (
            .O(N__43366),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__9668 (
            .O(N__43363),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__9667 (
            .O(N__43360),
            .I(N__43357));
    LocalMux I__9666 (
            .O(N__43357),
            .I(N__43354));
    Span4Mux_v I__9665 (
            .O(N__43354),
            .I(N__43351));
    Sp12to4 I__9664 (
            .O(N__43351),
            .I(N__43348));
    Span12Mux_h I__9663 (
            .O(N__43348),
            .I(N__43345));
    Odrv12 I__9662 (
            .O(N__43345),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    CascadeMux I__9661 (
            .O(N__43342),
            .I(N__43336));
    CascadeMux I__9660 (
            .O(N__43341),
            .I(N__43332));
    CascadeMux I__9659 (
            .O(N__43340),
            .I(N__43328));
    InMux I__9658 (
            .O(N__43339),
            .I(N__43324));
    InMux I__9657 (
            .O(N__43336),
            .I(N__43311));
    InMux I__9656 (
            .O(N__43335),
            .I(N__43311));
    InMux I__9655 (
            .O(N__43332),
            .I(N__43311));
    InMux I__9654 (
            .O(N__43331),
            .I(N__43311));
    InMux I__9653 (
            .O(N__43328),
            .I(N__43311));
    InMux I__9652 (
            .O(N__43327),
            .I(N__43311));
    LocalMux I__9651 (
            .O(N__43324),
            .I(N__43308));
    LocalMux I__9650 (
            .O(N__43311),
            .I(N__43304));
    Span12Mux_s7_v I__9649 (
            .O(N__43308),
            .I(N__43301));
    InMux I__9648 (
            .O(N__43307),
            .I(N__43298));
    Span4Mux_h I__9647 (
            .O(N__43304),
            .I(N__43295));
    Span12Mux_h I__9646 (
            .O(N__43301),
            .I(N__43290));
    LocalMux I__9645 (
            .O(N__43298),
            .I(N__43290));
    Span4Mux_h I__9644 (
            .O(N__43295),
            .I(N__43287));
    Span12Mux_h I__9643 (
            .O(N__43290),
            .I(N__43284));
    Span4Mux_h I__9642 (
            .O(N__43287),
            .I(N__43281));
    Odrv12 I__9641 (
            .O(N__43284),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    Odrv4 I__9640 (
            .O(N__43281),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    InMux I__9639 (
            .O(N__43276),
            .I(N__43273));
    LocalMux I__9638 (
            .O(N__43273),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__9637 (
            .O(N__43270),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__9636 (
            .O(N__43267),
            .I(N__43264));
    LocalMux I__9635 (
            .O(N__43264),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__9634 (
            .O(N__43261),
            .I(N__43258));
    LocalMux I__9633 (
            .O(N__43258),
            .I(N__43255));
    Span4Mux_v I__9632 (
            .O(N__43255),
            .I(N__43252));
    Odrv4 I__9631 (
            .O(N__43252),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__9630 (
            .O(N__43249),
            .I(bfn_16_29_0_));
    InMux I__9629 (
            .O(N__43246),
            .I(N__43243));
    LocalMux I__9628 (
            .O(N__43243),
            .I(N__43239));
    InMux I__9627 (
            .O(N__43242),
            .I(N__43236));
    Odrv4 I__9626 (
            .O(N__43239),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__9625 (
            .O(N__43236),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__9624 (
            .O(N__43231),
            .I(N__43228));
    LocalMux I__9623 (
            .O(N__43228),
            .I(N__43225));
    Span4Mux_v I__9622 (
            .O(N__43225),
            .I(N__43222));
    Odrv4 I__9621 (
            .O(N__43222),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__9620 (
            .O(N__43219),
            .I(N__43216));
    LocalMux I__9619 (
            .O(N__43216),
            .I(N__43213));
    Span4Mux_v I__9618 (
            .O(N__43213),
            .I(N__43210));
    Odrv4 I__9617 (
            .O(N__43210),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__9616 (
            .O(N__43207),
            .I(N__43202));
    InMux I__9615 (
            .O(N__43206),
            .I(N__43199));
    InMux I__9614 (
            .O(N__43205),
            .I(N__43196));
    LocalMux I__9613 (
            .O(N__43202),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__9612 (
            .O(N__43199),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__9611 (
            .O(N__43196),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__9610 (
            .O(N__43189),
            .I(N__43184));
    InMux I__9609 (
            .O(N__43188),
            .I(N__43181));
    InMux I__9608 (
            .O(N__43187),
            .I(N__43178));
    LocalMux I__9607 (
            .O(N__43184),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__9606 (
            .O(N__43181),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__9605 (
            .O(N__43178),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__9604 (
            .O(N__43171),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__9603 (
            .O(N__43168),
            .I(N__43165));
    LocalMux I__9602 (
            .O(N__43165),
            .I(N__43162));
    Span4Mux_v I__9601 (
            .O(N__43162),
            .I(N__43159));
    Sp12to4 I__9600 (
            .O(N__43159),
            .I(N__43156));
    Odrv12 I__9599 (
            .O(N__43156),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    CascadeMux I__9598 (
            .O(N__43153),
            .I(N__43150));
    InMux I__9597 (
            .O(N__43150),
            .I(N__43147));
    LocalMux I__9596 (
            .O(N__43147),
            .I(N__43144));
    Span4Mux_v I__9595 (
            .O(N__43144),
            .I(N__43141));
    Sp12to4 I__9594 (
            .O(N__43141),
            .I(N__43138));
    Span12Mux_h I__9593 (
            .O(N__43138),
            .I(N__43135));
    Odrv12 I__9592 (
            .O(N__43135),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    InMux I__9591 (
            .O(N__43132),
            .I(N__43129));
    LocalMux I__9590 (
            .O(N__43129),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__9589 (
            .O(N__43126),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__9588 (
            .O(N__43123),
            .I(N__43120));
    LocalMux I__9587 (
            .O(N__43120),
            .I(N__43117));
    Span4Mux_v I__9586 (
            .O(N__43117),
            .I(N__43114));
    Sp12to4 I__9585 (
            .O(N__43114),
            .I(N__43111));
    Odrv12 I__9584 (
            .O(N__43111),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    CascadeMux I__9583 (
            .O(N__43108),
            .I(N__43105));
    InMux I__9582 (
            .O(N__43105),
            .I(N__43102));
    LocalMux I__9581 (
            .O(N__43102),
            .I(N__43099));
    Span4Mux_v I__9580 (
            .O(N__43099),
            .I(N__43096));
    Span4Mux_h I__9579 (
            .O(N__43096),
            .I(N__43093));
    Span4Mux_h I__9578 (
            .O(N__43093),
            .I(N__43090));
    Span4Mux_h I__9577 (
            .O(N__43090),
            .I(N__43087));
    Odrv4 I__9576 (
            .O(N__43087),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__9575 (
            .O(N__43084),
            .I(N__43081));
    LocalMux I__9574 (
            .O(N__43081),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__9573 (
            .O(N__43078),
            .I(bfn_16_28_0_));
    InMux I__9572 (
            .O(N__43075),
            .I(N__43072));
    LocalMux I__9571 (
            .O(N__43072),
            .I(N__43069));
    Span4Mux_h I__9570 (
            .O(N__43069),
            .I(N__43066));
    Span4Mux_h I__9569 (
            .O(N__43066),
            .I(N__43063));
    Span4Mux_h I__9568 (
            .O(N__43063),
            .I(N__43060));
    Odrv4 I__9567 (
            .O(N__43060),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    CascadeMux I__9566 (
            .O(N__43057),
            .I(N__43054));
    InMux I__9565 (
            .O(N__43054),
            .I(N__43051));
    LocalMux I__9564 (
            .O(N__43051),
            .I(N__43048));
    Span4Mux_v I__9563 (
            .O(N__43048),
            .I(N__43045));
    Sp12to4 I__9562 (
            .O(N__43045),
            .I(N__43042));
    Span12Mux_h I__9561 (
            .O(N__43042),
            .I(N__43039));
    Odrv12 I__9560 (
            .O(N__43039),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__9559 (
            .O(N__43036),
            .I(N__43033));
    LocalMux I__9558 (
            .O(N__43033),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__9557 (
            .O(N__43030),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__9556 (
            .O(N__43027),
            .I(N__43024));
    InMux I__9555 (
            .O(N__43024),
            .I(N__43021));
    LocalMux I__9554 (
            .O(N__43021),
            .I(N__43018));
    Span4Mux_v I__9553 (
            .O(N__43018),
            .I(N__43015));
    Span4Mux_h I__9552 (
            .O(N__43015),
            .I(N__43012));
    Span4Mux_h I__9551 (
            .O(N__43012),
            .I(N__43009));
    Span4Mux_h I__9550 (
            .O(N__43009),
            .I(N__43006));
    Odrv4 I__9549 (
            .O(N__43006),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__9548 (
            .O(N__43003),
            .I(N__43000));
    LocalMux I__9547 (
            .O(N__43000),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__9546 (
            .O(N__42997),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__9545 (
            .O(N__42994),
            .I(N__42991));
    LocalMux I__9544 (
            .O(N__42991),
            .I(N__42988));
    Span4Mux_v I__9543 (
            .O(N__42988),
            .I(N__42985));
    Sp12to4 I__9542 (
            .O(N__42985),
            .I(N__42982));
    Span12Mux_h I__9541 (
            .O(N__42982),
            .I(N__42979));
    Odrv12 I__9540 (
            .O(N__42979),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__9539 (
            .O(N__42976),
            .I(N__42973));
    LocalMux I__9538 (
            .O(N__42973),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__9537 (
            .O(N__42970),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    CascadeMux I__9536 (
            .O(N__42967),
            .I(N__42964));
    InMux I__9535 (
            .O(N__42964),
            .I(N__42961));
    LocalMux I__9534 (
            .O(N__42961),
            .I(N__42958));
    Span12Mux_s6_v I__9533 (
            .O(N__42958),
            .I(N__42955));
    Span12Mux_h I__9532 (
            .O(N__42955),
            .I(N__42952));
    Odrv12 I__9531 (
            .O(N__42952),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__9530 (
            .O(N__42949),
            .I(N__42946));
    LocalMux I__9529 (
            .O(N__42946),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__9528 (
            .O(N__42943),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__9527 (
            .O(N__42940),
            .I(N__42937));
    LocalMux I__9526 (
            .O(N__42937),
            .I(N__42934));
    Span4Mux_h I__9525 (
            .O(N__42934),
            .I(N__42931));
    Span4Mux_v I__9524 (
            .O(N__42931),
            .I(N__42928));
    Sp12to4 I__9523 (
            .O(N__42928),
            .I(N__42925));
    Odrv12 I__9522 (
            .O(N__42925),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__9521 (
            .O(N__42922),
            .I(N__42919));
    LocalMux I__9520 (
            .O(N__42919),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__9519 (
            .O(N__42916),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__9518 (
            .O(N__42913),
            .I(N__42910));
    InMux I__9517 (
            .O(N__42910),
            .I(N__42906));
    InMux I__9516 (
            .O(N__42909),
            .I(N__42903));
    LocalMux I__9515 (
            .O(N__42906),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    LocalMux I__9514 (
            .O(N__42903),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__9513 (
            .O(N__42898),
            .I(N__42895));
    LocalMux I__9512 (
            .O(N__42895),
            .I(N__42892));
    Span4Mux_v I__9511 (
            .O(N__42892),
            .I(N__42889));
    Span4Mux_h I__9510 (
            .O(N__42889),
            .I(N__42886));
    Span4Mux_h I__9509 (
            .O(N__42886),
            .I(N__42883));
    Span4Mux_h I__9508 (
            .O(N__42883),
            .I(N__42880));
    Odrv4 I__9507 (
            .O(N__42880),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__9506 (
            .O(N__42877),
            .I(N__42874));
    InMux I__9505 (
            .O(N__42874),
            .I(N__42871));
    LocalMux I__9504 (
            .O(N__42871),
            .I(N__42868));
    Span4Mux_h I__9503 (
            .O(N__42868),
            .I(N__42865));
    Span4Mux_h I__9502 (
            .O(N__42865),
            .I(N__42862));
    Span4Mux_h I__9501 (
            .O(N__42862),
            .I(N__42859));
    Odrv4 I__9500 (
            .O(N__42859),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__9499 (
            .O(N__42856),
            .I(N__42853));
    LocalMux I__9498 (
            .O(N__42853),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__9497 (
            .O(N__42850),
            .I(N__42847));
    LocalMux I__9496 (
            .O(N__42847),
            .I(N__42844));
    Span4Mux_h I__9495 (
            .O(N__42844),
            .I(N__42841));
    Span4Mux_h I__9494 (
            .O(N__42841),
            .I(N__42838));
    Span4Mux_h I__9493 (
            .O(N__42838),
            .I(N__42835));
    Odrv4 I__9492 (
            .O(N__42835),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__9491 (
            .O(N__42832),
            .I(N__42829));
    InMux I__9490 (
            .O(N__42829),
            .I(N__42826));
    LocalMux I__9489 (
            .O(N__42826),
            .I(N__42823));
    Span4Mux_v I__9488 (
            .O(N__42823),
            .I(N__42820));
    Sp12to4 I__9487 (
            .O(N__42820),
            .I(N__42817));
    Span12Mux_h I__9486 (
            .O(N__42817),
            .I(N__42814));
    Odrv12 I__9485 (
            .O(N__42814),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__9484 (
            .O(N__42811),
            .I(N__42808));
    InMux I__9483 (
            .O(N__42808),
            .I(N__42805));
    LocalMux I__9482 (
            .O(N__42805),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__9481 (
            .O(N__42802),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__9480 (
            .O(N__42799),
            .I(N__42796));
    LocalMux I__9479 (
            .O(N__42796),
            .I(N__42793));
    Span4Mux_v I__9478 (
            .O(N__42793),
            .I(N__42790));
    Sp12to4 I__9477 (
            .O(N__42790),
            .I(N__42787));
    Span12Mux_h I__9476 (
            .O(N__42787),
            .I(N__42784));
    Odrv12 I__9475 (
            .O(N__42784),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__9474 (
            .O(N__42781),
            .I(N__42778));
    InMux I__9473 (
            .O(N__42778),
            .I(N__42775));
    LocalMux I__9472 (
            .O(N__42775),
            .I(N__42772));
    Span4Mux_h I__9471 (
            .O(N__42772),
            .I(N__42769));
    Span4Mux_h I__9470 (
            .O(N__42769),
            .I(N__42766));
    Span4Mux_h I__9469 (
            .O(N__42766),
            .I(N__42763));
    Odrv4 I__9468 (
            .O(N__42763),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__9467 (
            .O(N__42760),
            .I(N__42757));
    LocalMux I__9466 (
            .O(N__42757),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__9465 (
            .O(N__42754),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__9464 (
            .O(N__42751),
            .I(N__42748));
    LocalMux I__9463 (
            .O(N__42748),
            .I(N__42745));
    Span4Mux_v I__9462 (
            .O(N__42745),
            .I(N__42742));
    Sp12to4 I__9461 (
            .O(N__42742),
            .I(N__42739));
    Span12Mux_h I__9460 (
            .O(N__42739),
            .I(N__42736));
    Odrv12 I__9459 (
            .O(N__42736),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__9458 (
            .O(N__42733),
            .I(N__42730));
    InMux I__9457 (
            .O(N__42730),
            .I(N__42727));
    LocalMux I__9456 (
            .O(N__42727),
            .I(N__42724));
    Span12Mux_h I__9455 (
            .O(N__42724),
            .I(N__42721));
    Odrv12 I__9454 (
            .O(N__42721),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__9453 (
            .O(N__42718),
            .I(N__42715));
    InMux I__9452 (
            .O(N__42715),
            .I(N__42712));
    LocalMux I__9451 (
            .O(N__42712),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__9450 (
            .O(N__42709),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__9449 (
            .O(N__42706),
            .I(N__42703));
    LocalMux I__9448 (
            .O(N__42703),
            .I(N__42700));
    Span12Mux_s7_v I__9447 (
            .O(N__42700),
            .I(N__42697));
    Span12Mux_h I__9446 (
            .O(N__42697),
            .I(N__42694));
    Odrv12 I__9445 (
            .O(N__42694),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__9444 (
            .O(N__42691),
            .I(N__42688));
    InMux I__9443 (
            .O(N__42688),
            .I(N__42685));
    LocalMux I__9442 (
            .O(N__42685),
            .I(N__42682));
    Span4Mux_v I__9441 (
            .O(N__42682),
            .I(N__42679));
    Span4Mux_h I__9440 (
            .O(N__42679),
            .I(N__42676));
    Span4Mux_h I__9439 (
            .O(N__42676),
            .I(N__42673));
    Odrv4 I__9438 (
            .O(N__42673),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__9437 (
            .O(N__42670),
            .I(N__42667));
    LocalMux I__9436 (
            .O(N__42667),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__9435 (
            .O(N__42664),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__9434 (
            .O(N__42661),
            .I(N__42658));
    LocalMux I__9433 (
            .O(N__42658),
            .I(N__42655));
    Span4Mux_h I__9432 (
            .O(N__42655),
            .I(N__42652));
    Span4Mux_v I__9431 (
            .O(N__42652),
            .I(N__42649));
    Sp12to4 I__9430 (
            .O(N__42649),
            .I(N__42646));
    Odrv12 I__9429 (
            .O(N__42646),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__9428 (
            .O(N__42643),
            .I(N__42640));
    InMux I__9427 (
            .O(N__42640),
            .I(N__42637));
    LocalMux I__9426 (
            .O(N__42637),
            .I(N__42634));
    Span4Mux_v I__9425 (
            .O(N__42634),
            .I(N__42631));
    Sp12to4 I__9424 (
            .O(N__42631),
            .I(N__42628));
    Odrv12 I__9423 (
            .O(N__42628),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__9422 (
            .O(N__42625),
            .I(N__42622));
    LocalMux I__9421 (
            .O(N__42622),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__9420 (
            .O(N__42619),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__9419 (
            .O(N__42616),
            .I(N__42613));
    LocalMux I__9418 (
            .O(N__42613),
            .I(N__42610));
    Span12Mux_s5_v I__9417 (
            .O(N__42610),
            .I(N__42607));
    Odrv12 I__9416 (
            .O(N__42607),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    CascadeMux I__9415 (
            .O(N__42604),
            .I(N__42601));
    InMux I__9414 (
            .O(N__42601),
            .I(N__42598));
    LocalMux I__9413 (
            .O(N__42598),
            .I(N__42595));
    Span4Mux_v I__9412 (
            .O(N__42595),
            .I(N__42592));
    Sp12to4 I__9411 (
            .O(N__42592),
            .I(N__42589));
    Span12Mux_h I__9410 (
            .O(N__42589),
            .I(N__42586));
    Odrv12 I__9409 (
            .O(N__42586),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    InMux I__9408 (
            .O(N__42583),
            .I(N__42580));
    LocalMux I__9407 (
            .O(N__42580),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__9406 (
            .O(N__42577),
            .I(N__42574));
    LocalMux I__9405 (
            .O(N__42574),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__9404 (
            .O(N__42571),
            .I(N__42568));
    LocalMux I__9403 (
            .O(N__42568),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__9402 (
            .O(N__42565),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ));
    InMux I__9401 (
            .O(N__42562),
            .I(N__42559));
    LocalMux I__9400 (
            .O(N__42559),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__9399 (
            .O(N__42556),
            .I(N__42551));
    InMux I__9398 (
            .O(N__42555),
            .I(N__42548));
    InMux I__9397 (
            .O(N__42554),
            .I(N__42545));
    LocalMux I__9396 (
            .O(N__42551),
            .I(N__42538));
    LocalMux I__9395 (
            .O(N__42548),
            .I(N__42538));
    LocalMux I__9394 (
            .O(N__42545),
            .I(N__42538));
    Span4Mux_v I__9393 (
            .O(N__42538),
            .I(N__42535));
    Sp12to4 I__9392 (
            .O(N__42535),
            .I(N__42532));
    Span12Mux_h I__9391 (
            .O(N__42532),
            .I(N__42529));
    Span12Mux_v I__9390 (
            .O(N__42529),
            .I(N__42526));
    Odrv12 I__9389 (
            .O(N__42526),
            .I(il_min_comp2_c));
    InMux I__9388 (
            .O(N__42523),
            .I(N__42520));
    LocalMux I__9387 (
            .O(N__42520),
            .I(N__42517));
    Span4Mux_v I__9386 (
            .O(N__42517),
            .I(N__42513));
    InMux I__9385 (
            .O(N__42516),
            .I(N__42510));
    Span4Mux_v I__9384 (
            .O(N__42513),
            .I(N__42505));
    LocalMux I__9383 (
            .O(N__42510),
            .I(N__42505));
    Odrv4 I__9382 (
            .O(N__42505),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__9381 (
            .O(N__42502),
            .I(N__42498));
    CascadeMux I__9380 (
            .O(N__42501),
            .I(N__42495));
    LocalMux I__9379 (
            .O(N__42498),
            .I(N__42492));
    InMux I__9378 (
            .O(N__42495),
            .I(N__42488));
    Span4Mux_h I__9377 (
            .O(N__42492),
            .I(N__42485));
    InMux I__9376 (
            .O(N__42491),
            .I(N__42481));
    LocalMux I__9375 (
            .O(N__42488),
            .I(N__42478));
    Span4Mux_v I__9374 (
            .O(N__42485),
            .I(N__42475));
    InMux I__9373 (
            .O(N__42484),
            .I(N__42472));
    LocalMux I__9372 (
            .O(N__42481),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__9371 (
            .O(N__42478),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__9370 (
            .O(N__42475),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__9369 (
            .O(N__42472),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__9368 (
            .O(N__42463),
            .I(N__42458));
    InMux I__9367 (
            .O(N__42462),
            .I(N__42455));
    InMux I__9366 (
            .O(N__42461),
            .I(N__42452));
    LocalMux I__9365 (
            .O(N__42458),
            .I(N__42449));
    LocalMux I__9364 (
            .O(N__42455),
            .I(N__42444));
    LocalMux I__9363 (
            .O(N__42452),
            .I(N__42444));
    Span4Mux_v I__9362 (
            .O(N__42449),
            .I(N__42440));
    Span4Mux_v I__9361 (
            .O(N__42444),
            .I(N__42437));
    InMux I__9360 (
            .O(N__42443),
            .I(N__42432));
    Sp12to4 I__9359 (
            .O(N__42440),
            .I(N__42427));
    Sp12to4 I__9358 (
            .O(N__42437),
            .I(N__42427));
    InMux I__9357 (
            .O(N__42436),
            .I(N__42424));
    InMux I__9356 (
            .O(N__42435),
            .I(N__42420));
    LocalMux I__9355 (
            .O(N__42432),
            .I(N__42417));
    Span12Mux_h I__9354 (
            .O(N__42427),
            .I(N__42412));
    LocalMux I__9353 (
            .O(N__42424),
            .I(N__42412));
    InMux I__9352 (
            .O(N__42423),
            .I(N__42409));
    LocalMux I__9351 (
            .O(N__42420),
            .I(state_3));
    Odrv4 I__9350 (
            .O(N__42417),
            .I(state_3));
    Odrv12 I__9349 (
            .O(N__42412),
            .I(state_3));
    LocalMux I__9348 (
            .O(N__42409),
            .I(state_3));
    IoInMux I__9347 (
            .O(N__42400),
            .I(N__42397));
    LocalMux I__9346 (
            .O(N__42397),
            .I(N__42394));
    Span4Mux_s1_v I__9345 (
            .O(N__42394),
            .I(N__42391));
    Span4Mux_v I__9344 (
            .O(N__42391),
            .I(N__42388));
    Span4Mux_v I__9343 (
            .O(N__42388),
            .I(N__42384));
    InMux I__9342 (
            .O(N__42387),
            .I(N__42381));
    Odrv4 I__9341 (
            .O(N__42384),
            .I(test22_c));
    LocalMux I__9340 (
            .O(N__42381),
            .I(test22_c));
    InMux I__9339 (
            .O(N__42376),
            .I(N__42348));
    InMux I__9338 (
            .O(N__42375),
            .I(N__42331));
    InMux I__9337 (
            .O(N__42374),
            .I(N__42331));
    InMux I__9336 (
            .O(N__42373),
            .I(N__42331));
    InMux I__9335 (
            .O(N__42372),
            .I(N__42331));
    InMux I__9334 (
            .O(N__42371),
            .I(N__42331));
    InMux I__9333 (
            .O(N__42370),
            .I(N__42331));
    InMux I__9332 (
            .O(N__42369),
            .I(N__42331));
    InMux I__9331 (
            .O(N__42368),
            .I(N__42331));
    InMux I__9330 (
            .O(N__42367),
            .I(N__42316));
    InMux I__9329 (
            .O(N__42366),
            .I(N__42316));
    InMux I__9328 (
            .O(N__42365),
            .I(N__42316));
    InMux I__9327 (
            .O(N__42364),
            .I(N__42316));
    InMux I__9326 (
            .O(N__42363),
            .I(N__42316));
    InMux I__9325 (
            .O(N__42362),
            .I(N__42316));
    InMux I__9324 (
            .O(N__42361),
            .I(N__42316));
    CascadeMux I__9323 (
            .O(N__42360),
            .I(N__42313));
    CascadeMux I__9322 (
            .O(N__42359),
            .I(N__42306));
    CascadeMux I__9321 (
            .O(N__42358),
            .I(N__42302));
    CascadeMux I__9320 (
            .O(N__42357),
            .I(N__42299));
    CascadeMux I__9319 (
            .O(N__42356),
            .I(N__42296));
    InMux I__9318 (
            .O(N__42355),
            .I(N__42291));
    InMux I__9317 (
            .O(N__42354),
            .I(N__42291));
    InMux I__9316 (
            .O(N__42353),
            .I(N__42284));
    InMux I__9315 (
            .O(N__42352),
            .I(N__42284));
    InMux I__9314 (
            .O(N__42351),
            .I(N__42284));
    LocalMux I__9313 (
            .O(N__42348),
            .I(N__42277));
    LocalMux I__9312 (
            .O(N__42331),
            .I(N__42277));
    LocalMux I__9311 (
            .O(N__42316),
            .I(N__42277));
    InMux I__9310 (
            .O(N__42313),
            .I(N__42274));
    InMux I__9309 (
            .O(N__42312),
            .I(N__42271));
    InMux I__9308 (
            .O(N__42311),
            .I(N__42256));
    InMux I__9307 (
            .O(N__42310),
            .I(N__42256));
    InMux I__9306 (
            .O(N__42309),
            .I(N__42256));
    InMux I__9305 (
            .O(N__42306),
            .I(N__42256));
    InMux I__9304 (
            .O(N__42305),
            .I(N__42256));
    InMux I__9303 (
            .O(N__42302),
            .I(N__42256));
    InMux I__9302 (
            .O(N__42299),
            .I(N__42256));
    InMux I__9301 (
            .O(N__42296),
            .I(N__42253));
    LocalMux I__9300 (
            .O(N__42291),
            .I(N__42247));
    LocalMux I__9299 (
            .O(N__42284),
            .I(N__42247));
    Span4Mux_v I__9298 (
            .O(N__42277),
            .I(N__42244));
    LocalMux I__9297 (
            .O(N__42274),
            .I(N__42239));
    LocalMux I__9296 (
            .O(N__42271),
            .I(N__42239));
    LocalMux I__9295 (
            .O(N__42256),
            .I(N__42236));
    LocalMux I__9294 (
            .O(N__42253),
            .I(N__42233));
    CascadeMux I__9293 (
            .O(N__42252),
            .I(N__42230));
    Span4Mux_v I__9292 (
            .O(N__42247),
            .I(N__42227));
    Sp12to4 I__9291 (
            .O(N__42244),
            .I(N__42224));
    Span4Mux_v I__9290 (
            .O(N__42239),
            .I(N__42221));
    Span4Mux_h I__9289 (
            .O(N__42236),
            .I(N__42218));
    Span4Mux_h I__9288 (
            .O(N__42233),
            .I(N__42215));
    InMux I__9287 (
            .O(N__42230),
            .I(N__42212));
    Sp12to4 I__9286 (
            .O(N__42227),
            .I(N__42209));
    Span12Mux_s8_h I__9285 (
            .O(N__42224),
            .I(N__42206));
    Odrv4 I__9284 (
            .O(N__42221),
            .I(N_19_1));
    Odrv4 I__9283 (
            .O(N__42218),
            .I(N_19_1));
    Odrv4 I__9282 (
            .O(N__42215),
            .I(N_19_1));
    LocalMux I__9281 (
            .O(N__42212),
            .I(N_19_1));
    Odrv12 I__9280 (
            .O(N__42209),
            .I(N_19_1));
    Odrv12 I__9279 (
            .O(N__42206),
            .I(N_19_1));
    InMux I__9278 (
            .O(N__42193),
            .I(N__42189));
    InMux I__9277 (
            .O(N__42192),
            .I(N__42186));
    LocalMux I__9276 (
            .O(N__42189),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    LocalMux I__9275 (
            .O(N__42186),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__9274 (
            .O(N__42181),
            .I(N__42175));
    InMux I__9273 (
            .O(N__42180),
            .I(N__42175));
    LocalMux I__9272 (
            .O(N__42175),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    CascadeMux I__9271 (
            .O(N__42172),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ));
    InMux I__9270 (
            .O(N__42169),
            .I(N__42166));
    LocalMux I__9269 (
            .O(N__42166),
            .I(N__42163));
    Odrv12 I__9268 (
            .O(N__42163),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__9267 (
            .O(N__42160),
            .I(N__42156));
    InMux I__9266 (
            .O(N__42159),
            .I(N__42153));
    LocalMux I__9265 (
            .O(N__42156),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__9264 (
            .O(N__42153),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__9263 (
            .O(N__42148),
            .I(N__42141));
    InMux I__9262 (
            .O(N__42147),
            .I(N__42141));
    InMux I__9261 (
            .O(N__42146),
            .I(N__42137));
    LocalMux I__9260 (
            .O(N__42141),
            .I(N__42134));
    InMux I__9259 (
            .O(N__42140),
            .I(N__42131));
    LocalMux I__9258 (
            .O(N__42137),
            .I(N__42128));
    Span4Mux_h I__9257 (
            .O(N__42134),
            .I(N__42125));
    LocalMux I__9256 (
            .O(N__42131),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv12 I__9255 (
            .O(N__42128),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__9254 (
            .O(N__42125),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__9253 (
            .O(N__42118),
            .I(N__42115));
    InMux I__9252 (
            .O(N__42115),
            .I(N__42112));
    LocalMux I__9251 (
            .O(N__42112),
            .I(N__42108));
    InMux I__9250 (
            .O(N__42111),
            .I(N__42105));
    Odrv4 I__9249 (
            .O(N__42108),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    LocalMux I__9248 (
            .O(N__42105),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__9247 (
            .O(N__42100),
            .I(N__42097));
    LocalMux I__9246 (
            .O(N__42097),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    CascadeMux I__9245 (
            .O(N__42094),
            .I(N__42090));
    InMux I__9244 (
            .O(N__42093),
            .I(N__42087));
    InMux I__9243 (
            .O(N__42090),
            .I(N__42082));
    LocalMux I__9242 (
            .O(N__42087),
            .I(N__42079));
    InMux I__9241 (
            .O(N__42086),
            .I(N__42074));
    InMux I__9240 (
            .O(N__42085),
            .I(N__42074));
    LocalMux I__9239 (
            .O(N__42082),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__9238 (
            .O(N__42079),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__9237 (
            .O(N__42074),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__9236 (
            .O(N__42067),
            .I(N__42064));
    InMux I__9235 (
            .O(N__42064),
            .I(N__42061));
    LocalMux I__9234 (
            .O(N__42061),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    InMux I__9233 (
            .O(N__42058),
            .I(N__42055));
    LocalMux I__9232 (
            .O(N__42055),
            .I(N__42052));
    Span4Mux_h I__9231 (
            .O(N__42052),
            .I(N__42049));
    Odrv4 I__9230 (
            .O(N__42049),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0 ));
    InMux I__9229 (
            .O(N__42046),
            .I(N__42042));
    InMux I__9228 (
            .O(N__42045),
            .I(N__42039));
    LocalMux I__9227 (
            .O(N__42042),
            .I(N__42034));
    LocalMux I__9226 (
            .O(N__42039),
            .I(N__42034));
    Span4Mux_v I__9225 (
            .O(N__42034),
            .I(N__42030));
    InMux I__9224 (
            .O(N__42033),
            .I(N__42027));
    Sp12to4 I__9223 (
            .O(N__42030),
            .I(N__42022));
    LocalMux I__9222 (
            .O(N__42027),
            .I(N__42022));
    Span12Mux_h I__9221 (
            .O(N__42022),
            .I(N__42019));
    Span12Mux_v I__9220 (
            .O(N__42019),
            .I(N__42016));
    Odrv12 I__9219 (
            .O(N__42016),
            .I(il_max_comp2_c));
    InMux I__9218 (
            .O(N__42013),
            .I(N__42010));
    LocalMux I__9217 (
            .O(N__42010),
            .I(N__42006));
    CascadeMux I__9216 (
            .O(N__42009),
            .I(N__42002));
    Span4Mux_v I__9215 (
            .O(N__42006),
            .I(N__41999));
    CascadeMux I__9214 (
            .O(N__42005),
            .I(N__41996));
    InMux I__9213 (
            .O(N__42002),
            .I(N__41993));
    Span4Mux_h I__9212 (
            .O(N__41999),
            .I(N__41990));
    InMux I__9211 (
            .O(N__41996),
            .I(N__41986));
    LocalMux I__9210 (
            .O(N__41993),
            .I(N__41981));
    Span4Mux_v I__9209 (
            .O(N__41990),
            .I(N__41981));
    InMux I__9208 (
            .O(N__41989),
            .I(N__41978));
    LocalMux I__9207 (
            .O(N__41986),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__9206 (
            .O(N__41981),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__9205 (
            .O(N__41978),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__9204 (
            .O(N__41971),
            .I(N__41968));
    LocalMux I__9203 (
            .O(N__41968),
            .I(N__41964));
    InMux I__9202 (
            .O(N__41967),
            .I(N__41961));
    Span4Mux_h I__9201 (
            .O(N__41964),
            .I(N__41958));
    LocalMux I__9200 (
            .O(N__41961),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    Odrv4 I__9199 (
            .O(N__41958),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__9198 (
            .O(N__41953),
            .I(N__41950));
    LocalMux I__9197 (
            .O(N__41950),
            .I(N__41946));
    InMux I__9196 (
            .O(N__41949),
            .I(N__41943));
    Odrv4 I__9195 (
            .O(N__41946),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__9194 (
            .O(N__41943),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__9193 (
            .O(N__41938),
            .I(N__41935));
    InMux I__9192 (
            .O(N__41935),
            .I(N__41932));
    LocalMux I__9191 (
            .O(N__41932),
            .I(N__41928));
    InMux I__9190 (
            .O(N__41931),
            .I(N__41925));
    Odrv4 I__9189 (
            .O(N__41928),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__9188 (
            .O(N__41925),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__9187 (
            .O(N__41920),
            .I(N__41917));
    LocalMux I__9186 (
            .O(N__41917),
            .I(N__41914));
    Span4Mux_h I__9185 (
            .O(N__41914),
            .I(N__41910));
    InMux I__9184 (
            .O(N__41913),
            .I(N__41907));
    Odrv4 I__9183 (
            .O(N__41910),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__9182 (
            .O(N__41907),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__9181 (
            .O(N__41902),
            .I(N__41899));
    LocalMux I__9180 (
            .O(N__41899),
            .I(N__41895));
    InMux I__9179 (
            .O(N__41898),
            .I(N__41892));
    Span4Mux_v I__9178 (
            .O(N__41895),
            .I(N__41889));
    LocalMux I__9177 (
            .O(N__41892),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__9176 (
            .O(N__41889),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__9175 (
            .O(N__41884),
            .I(N__41881));
    LocalMux I__9174 (
            .O(N__41881),
            .I(N__41875));
    InMux I__9173 (
            .O(N__41880),
            .I(N__41870));
    InMux I__9172 (
            .O(N__41879),
            .I(N__41870));
    InMux I__9171 (
            .O(N__41878),
            .I(N__41867));
    Span4Mux_h I__9170 (
            .O(N__41875),
            .I(N__41862));
    LocalMux I__9169 (
            .O(N__41870),
            .I(N__41862));
    LocalMux I__9168 (
            .O(N__41867),
            .I(N__41859));
    Odrv4 I__9167 (
            .O(N__41862),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__9166 (
            .O(N__41859),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    CascadeMux I__9165 (
            .O(N__41854),
            .I(N__41851));
    InMux I__9164 (
            .O(N__41851),
            .I(N__41845));
    InMux I__9163 (
            .O(N__41850),
            .I(N__41845));
    LocalMux I__9162 (
            .O(N__41845),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__9161 (
            .O(N__41842),
            .I(N__41838));
    InMux I__9160 (
            .O(N__41841),
            .I(N__41835));
    LocalMux I__9159 (
            .O(N__41838),
            .I(N__41831));
    LocalMux I__9158 (
            .O(N__41835),
            .I(N__41828));
    InMux I__9157 (
            .O(N__41834),
            .I(N__41825));
    Odrv12 I__9156 (
            .O(N__41831),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__9155 (
            .O(N__41828),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    LocalMux I__9154 (
            .O(N__41825),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__9153 (
            .O(N__41818),
            .I(N__41815));
    InMux I__9152 (
            .O(N__41815),
            .I(N__41811));
    InMux I__9151 (
            .O(N__41814),
            .I(N__41808));
    LocalMux I__9150 (
            .O(N__41811),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__9149 (
            .O(N__41808),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    CascadeMux I__9148 (
            .O(N__41803),
            .I(N__41798));
    InMux I__9147 (
            .O(N__41802),
            .I(N__41795));
    InMux I__9146 (
            .O(N__41801),
            .I(N__41790));
    InMux I__9145 (
            .O(N__41798),
            .I(N__41787));
    LocalMux I__9144 (
            .O(N__41795),
            .I(N__41784));
    InMux I__9143 (
            .O(N__41794),
            .I(N__41779));
    InMux I__9142 (
            .O(N__41793),
            .I(N__41779));
    LocalMux I__9141 (
            .O(N__41790),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__9140 (
            .O(N__41787),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__9139 (
            .O(N__41784),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__9138 (
            .O(N__41779),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__9137 (
            .O(N__41770),
            .I(N__41767));
    LocalMux I__9136 (
            .O(N__41767),
            .I(N__41762));
    InMux I__9135 (
            .O(N__41766),
            .I(N__41755));
    InMux I__9134 (
            .O(N__41765),
            .I(N__41755));
    Span4Mux_h I__9133 (
            .O(N__41762),
            .I(N__41752));
    InMux I__9132 (
            .O(N__41761),
            .I(N__41749));
    InMux I__9131 (
            .O(N__41760),
            .I(N__41746));
    LocalMux I__9130 (
            .O(N__41755),
            .I(N__41743));
    Odrv4 I__9129 (
            .O(N__41752),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__9128 (
            .O(N__41749),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__9127 (
            .O(N__41746),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__9126 (
            .O(N__41743),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__9125 (
            .O(N__41734),
            .I(N__41731));
    LocalMux I__9124 (
            .O(N__41731),
            .I(N__41727));
    InMux I__9123 (
            .O(N__41730),
            .I(N__41724));
    Odrv4 I__9122 (
            .O(N__41727),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    LocalMux I__9121 (
            .O(N__41724),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    InMux I__9120 (
            .O(N__41719),
            .I(N__41714));
    InMux I__9119 (
            .O(N__41718),
            .I(N__41711));
    InMux I__9118 (
            .O(N__41717),
            .I(N__41708));
    LocalMux I__9117 (
            .O(N__41714),
            .I(N__41705));
    LocalMux I__9116 (
            .O(N__41711),
            .I(N__41700));
    LocalMux I__9115 (
            .O(N__41708),
            .I(N__41700));
    Span4Mux_v I__9114 (
            .O(N__41705),
            .I(N__41697));
    Span4Mux_v I__9113 (
            .O(N__41700),
            .I(N__41694));
    Sp12to4 I__9112 (
            .O(N__41697),
            .I(N__41689));
    Sp12to4 I__9111 (
            .O(N__41694),
            .I(N__41689));
    Span12Mux_h I__9110 (
            .O(N__41689),
            .I(N__41686));
    Span12Mux_v I__9109 (
            .O(N__41686),
            .I(N__41683));
    Odrv12 I__9108 (
            .O(N__41683),
            .I(il_max_comp1_c));
    InMux I__9107 (
            .O(N__41680),
            .I(N__41673));
    InMux I__9106 (
            .O(N__41679),
            .I(N__41673));
    InMux I__9105 (
            .O(N__41678),
            .I(N__41670));
    LocalMux I__9104 (
            .O(N__41673),
            .I(N__41665));
    LocalMux I__9103 (
            .O(N__41670),
            .I(N__41665));
    Span4Mux_v I__9102 (
            .O(N__41665),
            .I(N__41662));
    Sp12to4 I__9101 (
            .O(N__41662),
            .I(N__41659));
    Span12Mux_h I__9100 (
            .O(N__41659),
            .I(N__41656));
    Span12Mux_v I__9099 (
            .O(N__41656),
            .I(N__41653));
    Odrv12 I__9098 (
            .O(N__41653),
            .I(il_min_comp1_c));
    CascadeMux I__9097 (
            .O(N__41650),
            .I(N__41647));
    InMux I__9096 (
            .O(N__41647),
            .I(N__41643));
    InMux I__9095 (
            .O(N__41646),
            .I(N__41639));
    LocalMux I__9094 (
            .O(N__41643),
            .I(N__41636));
    InMux I__9093 (
            .O(N__41642),
            .I(N__41633));
    LocalMux I__9092 (
            .O(N__41639),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__9091 (
            .O(N__41636),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__9090 (
            .O(N__41633),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__9089 (
            .O(N__41626),
            .I(N__41623));
    LocalMux I__9088 (
            .O(N__41623),
            .I(N__41620));
    Span4Mux_v I__9087 (
            .O(N__41620),
            .I(N__41614));
    InMux I__9086 (
            .O(N__41619),
            .I(N__41609));
    InMux I__9085 (
            .O(N__41618),
            .I(N__41609));
    InMux I__9084 (
            .O(N__41617),
            .I(N__41606));
    Odrv4 I__9083 (
            .O(N__41614),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__9082 (
            .O(N__41609),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__9081 (
            .O(N__41606),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__9080 (
            .O(N__41599),
            .I(N__41595));
    InMux I__9079 (
            .O(N__41598),
            .I(N__41592));
    LocalMux I__9078 (
            .O(N__41595),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__9077 (
            .O(N__41592),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__9076 (
            .O(N__41587),
            .I(N__41584));
    LocalMux I__9075 (
            .O(N__41584),
            .I(N__41579));
    InMux I__9074 (
            .O(N__41583),
            .I(N__41573));
    InMux I__9073 (
            .O(N__41582),
            .I(N__41573));
    Span4Mux_v I__9072 (
            .O(N__41579),
            .I(N__41570));
    InMux I__9071 (
            .O(N__41578),
            .I(N__41567));
    LocalMux I__9070 (
            .O(N__41573),
            .I(N__41564));
    Odrv4 I__9069 (
            .O(N__41570),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__9068 (
            .O(N__41567),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__9067 (
            .O(N__41564),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__9066 (
            .O(N__41557),
            .I(N__41554));
    LocalMux I__9065 (
            .O(N__41554),
            .I(N__41550));
    InMux I__9064 (
            .O(N__41553),
            .I(N__41547));
    Odrv4 I__9063 (
            .O(N__41550),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__9062 (
            .O(N__41547),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__9061 (
            .O(N__41542),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_ ));
    InMux I__9060 (
            .O(N__41539),
            .I(N__41534));
    InMux I__9059 (
            .O(N__41538),
            .I(N__41531));
    InMux I__9058 (
            .O(N__41537),
            .I(N__41528));
    LocalMux I__9057 (
            .O(N__41534),
            .I(N__41523));
    LocalMux I__9056 (
            .O(N__41531),
            .I(N__41523));
    LocalMux I__9055 (
            .O(N__41528),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv12 I__9054 (
            .O(N__41523),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__9053 (
            .O(N__41518),
            .I(N__41513));
    InMux I__9052 (
            .O(N__41517),
            .I(N__41510));
    InMux I__9051 (
            .O(N__41516),
            .I(N__41507));
    LocalMux I__9050 (
            .O(N__41513),
            .I(N__41504));
    LocalMux I__9049 (
            .O(N__41510),
            .I(N__41501));
    LocalMux I__9048 (
            .O(N__41507),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    Odrv4 I__9047 (
            .O(N__41504),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    Odrv4 I__9046 (
            .O(N__41501),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    InMux I__9045 (
            .O(N__41494),
            .I(N__41490));
    InMux I__9044 (
            .O(N__41493),
            .I(N__41486));
    LocalMux I__9043 (
            .O(N__41490),
            .I(N__41482));
    InMux I__9042 (
            .O(N__41489),
            .I(N__41479));
    LocalMux I__9041 (
            .O(N__41486),
            .I(N__41476));
    InMux I__9040 (
            .O(N__41485),
            .I(N__41473));
    Span4Mux_v I__9039 (
            .O(N__41482),
            .I(N__41470));
    LocalMux I__9038 (
            .O(N__41479),
            .I(N__41465));
    Span4Mux_h I__9037 (
            .O(N__41476),
            .I(N__41465));
    LocalMux I__9036 (
            .O(N__41473),
            .I(N__41462));
    Odrv4 I__9035 (
            .O(N__41470),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__9034 (
            .O(N__41465),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__9033 (
            .O(N__41462),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9032 (
            .O(N__41455),
            .I(N__41449));
    InMux I__9031 (
            .O(N__41454),
            .I(N__41449));
    LocalMux I__9030 (
            .O(N__41449),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    InMux I__9029 (
            .O(N__41446),
            .I(N__41441));
    InMux I__9028 (
            .O(N__41445),
            .I(N__41438));
    InMux I__9027 (
            .O(N__41444),
            .I(N__41435));
    LocalMux I__9026 (
            .O(N__41441),
            .I(N__41432));
    LocalMux I__9025 (
            .O(N__41438),
            .I(N__41428));
    LocalMux I__9024 (
            .O(N__41435),
            .I(N__41425));
    Span4Mux_v I__9023 (
            .O(N__41432),
            .I(N__41422));
    InMux I__9022 (
            .O(N__41431),
            .I(N__41419));
    Span4Mux_h I__9021 (
            .O(N__41428),
            .I(N__41414));
    Span4Mux_h I__9020 (
            .O(N__41425),
            .I(N__41414));
    Odrv4 I__9019 (
            .O(N__41422),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__9018 (
            .O(N__41419),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__9017 (
            .O(N__41414),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__9016 (
            .O(N__41407),
            .I(N__41402));
    InMux I__9015 (
            .O(N__41406),
            .I(N__41399));
    InMux I__9014 (
            .O(N__41405),
            .I(N__41396));
    LocalMux I__9013 (
            .O(N__41402),
            .I(N__41393));
    LocalMux I__9012 (
            .O(N__41399),
            .I(N__41390));
    LocalMux I__9011 (
            .O(N__41396),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv4 I__9010 (
            .O(N__41393),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv12 I__9009 (
            .O(N__41390),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__9008 (
            .O(N__41383),
            .I(N__41380));
    InMux I__9007 (
            .O(N__41380),
            .I(N__41374));
    InMux I__9006 (
            .O(N__41379),
            .I(N__41374));
    LocalMux I__9005 (
            .O(N__41374),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    InMux I__9004 (
            .O(N__41371),
            .I(N__41365));
    InMux I__9003 (
            .O(N__41370),
            .I(N__41365));
    LocalMux I__9002 (
            .O(N__41365),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__9001 (
            .O(N__41362),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__9000 (
            .O(N__41359),
            .I(N__41356));
    LocalMux I__8999 (
            .O(N__41356),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__8998 (
            .O(N__41353),
            .I(N__41347));
    InMux I__8997 (
            .O(N__41352),
            .I(N__41347));
    LocalMux I__8996 (
            .O(N__41347),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__8995 (
            .O(N__41344),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__8994 (
            .O(N__41341),
            .I(N__41338));
    LocalMux I__8993 (
            .O(N__41338),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__8992 (
            .O(N__41335),
            .I(N__41332));
    LocalMux I__8991 (
            .O(N__41332),
            .I(N__41329));
    Span4Mux_h I__8990 (
            .O(N__41329),
            .I(N__41325));
    InMux I__8989 (
            .O(N__41328),
            .I(N__41322));
    Odrv4 I__8988 (
            .O(N__41325),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__8987 (
            .O(N__41322),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__8986 (
            .O(N__41317),
            .I(N__41314));
    InMux I__8985 (
            .O(N__41314),
            .I(N__41311));
    LocalMux I__8984 (
            .O(N__41311),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ));
    InMux I__8983 (
            .O(N__41308),
            .I(N__41304));
    CascadeMux I__8982 (
            .O(N__41307),
            .I(N__41300));
    LocalMux I__8981 (
            .O(N__41304),
            .I(N__41297));
    InMux I__8980 (
            .O(N__41303),
            .I(N__41292));
    InMux I__8979 (
            .O(N__41300),
            .I(N__41289));
    Span4Mux_h I__8978 (
            .O(N__41297),
            .I(N__41286));
    InMux I__8977 (
            .O(N__41296),
            .I(N__41281));
    InMux I__8976 (
            .O(N__41295),
            .I(N__41281));
    LocalMux I__8975 (
            .O(N__41292),
            .I(N__41278));
    LocalMux I__8974 (
            .O(N__41289),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8973 (
            .O(N__41286),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__8972 (
            .O(N__41281),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8971 (
            .O(N__41278),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    IoInMux I__8970 (
            .O(N__41269),
            .I(N__41266));
    LocalMux I__8969 (
            .O(N__41266),
            .I(N__41263));
    Span4Mux_s1_v I__8968 (
            .O(N__41263),
            .I(N__41234));
    InMux I__8967 (
            .O(N__41262),
            .I(N__41223));
    InMux I__8966 (
            .O(N__41261),
            .I(N__41223));
    InMux I__8965 (
            .O(N__41260),
            .I(N__41223));
    InMux I__8964 (
            .O(N__41259),
            .I(N__41214));
    InMux I__8963 (
            .O(N__41258),
            .I(N__41214));
    InMux I__8962 (
            .O(N__41257),
            .I(N__41214));
    InMux I__8961 (
            .O(N__41256),
            .I(N__41214));
    InMux I__8960 (
            .O(N__41255),
            .I(N__41205));
    InMux I__8959 (
            .O(N__41254),
            .I(N__41205));
    InMux I__8958 (
            .O(N__41253),
            .I(N__41205));
    InMux I__8957 (
            .O(N__41252),
            .I(N__41205));
    InMux I__8956 (
            .O(N__41251),
            .I(N__41196));
    InMux I__8955 (
            .O(N__41250),
            .I(N__41196));
    InMux I__8954 (
            .O(N__41249),
            .I(N__41196));
    InMux I__8953 (
            .O(N__41248),
            .I(N__41196));
    InMux I__8952 (
            .O(N__41247),
            .I(N__41187));
    InMux I__8951 (
            .O(N__41246),
            .I(N__41187));
    InMux I__8950 (
            .O(N__41245),
            .I(N__41187));
    InMux I__8949 (
            .O(N__41244),
            .I(N__41187));
    InMux I__8948 (
            .O(N__41243),
            .I(N__41178));
    InMux I__8947 (
            .O(N__41242),
            .I(N__41178));
    InMux I__8946 (
            .O(N__41241),
            .I(N__41178));
    InMux I__8945 (
            .O(N__41240),
            .I(N__41178));
    InMux I__8944 (
            .O(N__41239),
            .I(N__41171));
    InMux I__8943 (
            .O(N__41238),
            .I(N__41171));
    InMux I__8942 (
            .O(N__41237),
            .I(N__41171));
    Span4Mux_v I__8941 (
            .O(N__41234),
            .I(N__41168));
    InMux I__8940 (
            .O(N__41233),
            .I(N__41159));
    InMux I__8939 (
            .O(N__41232),
            .I(N__41159));
    InMux I__8938 (
            .O(N__41231),
            .I(N__41159));
    InMux I__8937 (
            .O(N__41230),
            .I(N__41159));
    LocalMux I__8936 (
            .O(N__41223),
            .I(N__41156));
    LocalMux I__8935 (
            .O(N__41214),
            .I(N__41145));
    LocalMux I__8934 (
            .O(N__41205),
            .I(N__41145));
    LocalMux I__8933 (
            .O(N__41196),
            .I(N__41145));
    LocalMux I__8932 (
            .O(N__41187),
            .I(N__41145));
    LocalMux I__8931 (
            .O(N__41178),
            .I(N__41145));
    LocalMux I__8930 (
            .O(N__41171),
            .I(N__41142));
    Sp12to4 I__8929 (
            .O(N__41168),
            .I(N__41139));
    LocalMux I__8928 (
            .O(N__41159),
            .I(N__41130));
    Span4Mux_v I__8927 (
            .O(N__41156),
            .I(N__41130));
    Span4Mux_v I__8926 (
            .O(N__41145),
            .I(N__41130));
    Span4Mux_v I__8925 (
            .O(N__41142),
            .I(N__41130));
    Span12Mux_h I__8924 (
            .O(N__41139),
            .I(N__41127));
    Span4Mux_h I__8923 (
            .O(N__41130),
            .I(N__41124));
    Span12Mux_v I__8922 (
            .O(N__41127),
            .I(N__41121));
    Odrv4 I__8921 (
            .O(N__41124),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__8920 (
            .O(N__41121),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__8919 (
            .O(N__41116),
            .I(N__41113));
    LocalMux I__8918 (
            .O(N__41113),
            .I(N__41110));
    Sp12to4 I__8917 (
            .O(N__41110),
            .I(N__41107));
    Odrv12 I__8916 (
            .O(N__41107),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8915 (
            .O(N__41104),
            .I(N__41101));
    InMux I__8914 (
            .O(N__41101),
            .I(N__41098));
    LocalMux I__8913 (
            .O(N__41098),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__8912 (
            .O(N__41095),
            .I(N__41092));
    InMux I__8911 (
            .O(N__41092),
            .I(N__41089));
    LocalMux I__8910 (
            .O(N__41089),
            .I(N__41086));
    Odrv4 I__8909 (
            .O(N__41086),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__8908 (
            .O(N__41083),
            .I(N__41080));
    InMux I__8907 (
            .O(N__41080),
            .I(N__41077));
    LocalMux I__8906 (
            .O(N__41077),
            .I(N__41074));
    Span4Mux_h I__8905 (
            .O(N__41074),
            .I(N__41071));
    Odrv4 I__8904 (
            .O(N__41071),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    InMux I__8903 (
            .O(N__41068),
            .I(N__41062));
    InMux I__8902 (
            .O(N__41067),
            .I(N__41062));
    LocalMux I__8901 (
            .O(N__41062),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__8900 (
            .O(N__41059),
            .I(N__41055));
    InMux I__8899 (
            .O(N__41058),
            .I(N__41050));
    InMux I__8898 (
            .O(N__41055),
            .I(N__41050));
    LocalMux I__8897 (
            .O(N__41050),
            .I(N__41046));
    InMux I__8896 (
            .O(N__41049),
            .I(N__41043));
    Span4Mux_v I__8895 (
            .O(N__41046),
            .I(N__41040));
    LocalMux I__8894 (
            .O(N__41043),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__8893 (
            .O(N__41040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    CascadeMux I__8892 (
            .O(N__41035),
            .I(N__41032));
    InMux I__8891 (
            .O(N__41032),
            .I(N__41028));
    InMux I__8890 (
            .O(N__41031),
            .I(N__41025));
    LocalMux I__8889 (
            .O(N__41028),
            .I(N__41019));
    LocalMux I__8888 (
            .O(N__41025),
            .I(N__41019));
    InMux I__8887 (
            .O(N__41024),
            .I(N__41016));
    Span4Mux_v I__8886 (
            .O(N__41019),
            .I(N__41013));
    LocalMux I__8885 (
            .O(N__41016),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__8884 (
            .O(N__41013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__8883 (
            .O(N__41008),
            .I(N__41004));
    InMux I__8882 (
            .O(N__41007),
            .I(N__41001));
    LocalMux I__8881 (
            .O(N__41004),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    LocalMux I__8880 (
            .O(N__41001),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__8879 (
            .O(N__40996),
            .I(N__40993));
    LocalMux I__8878 (
            .O(N__40993),
            .I(N__40990));
    Odrv4 I__8877 (
            .O(N__40990),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    InMux I__8876 (
            .O(N__40987),
            .I(N__40984));
    LocalMux I__8875 (
            .O(N__40984),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__8874 (
            .O(N__40981),
            .I(N__40978));
    InMux I__8873 (
            .O(N__40978),
            .I(N__40975));
    LocalMux I__8872 (
            .O(N__40975),
            .I(N__40972));
    Odrv4 I__8871 (
            .O(N__40972),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__8870 (
            .O(N__40969),
            .I(N__40963));
    InMux I__8869 (
            .O(N__40968),
            .I(N__40963));
    LocalMux I__8868 (
            .O(N__40963),
            .I(N__40959));
    InMux I__8867 (
            .O(N__40962),
            .I(N__40956));
    Span4Mux_h I__8866 (
            .O(N__40959),
            .I(N__40953));
    LocalMux I__8865 (
            .O(N__40956),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__8864 (
            .O(N__40953),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__8863 (
            .O(N__40948),
            .I(N__40945));
    InMux I__8862 (
            .O(N__40945),
            .I(N__40939));
    InMux I__8861 (
            .O(N__40944),
            .I(N__40939));
    LocalMux I__8860 (
            .O(N__40939),
            .I(N__40935));
    InMux I__8859 (
            .O(N__40938),
            .I(N__40932));
    Span4Mux_h I__8858 (
            .O(N__40935),
            .I(N__40929));
    LocalMux I__8857 (
            .O(N__40932),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__8856 (
            .O(N__40929),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__8855 (
            .O(N__40924),
            .I(N__40921));
    InMux I__8854 (
            .O(N__40921),
            .I(N__40915));
    InMux I__8853 (
            .O(N__40920),
            .I(N__40915));
    LocalMux I__8852 (
            .O(N__40915),
            .I(N__40912));
    Odrv4 I__8851 (
            .O(N__40912),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8850 (
            .O(N__40909),
            .I(N__40906));
    LocalMux I__8849 (
            .O(N__40906),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__8848 (
            .O(N__40903),
            .I(N__40900));
    LocalMux I__8847 (
            .O(N__40900),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__8846 (
            .O(N__40897),
            .I(N__40894));
    LocalMux I__8845 (
            .O(N__40894),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    CascadeMux I__8844 (
            .O(N__40891),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ));
    InMux I__8843 (
            .O(N__40888),
            .I(N__40885));
    LocalMux I__8842 (
            .O(N__40885),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    InMux I__8841 (
            .O(N__40882),
            .I(N__40879));
    LocalMux I__8840 (
            .O(N__40879),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    CascadeMux I__8839 (
            .O(N__40876),
            .I(N__40873));
    InMux I__8838 (
            .O(N__40873),
            .I(N__40870));
    LocalMux I__8837 (
            .O(N__40870),
            .I(N__40867));
    Span4Mux_h I__8836 (
            .O(N__40867),
            .I(N__40864));
    Odrv4 I__8835 (
            .O(N__40864),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__8834 (
            .O(N__40861),
            .I(N__40857));
    InMux I__8833 (
            .O(N__40860),
            .I(N__40852));
    InMux I__8832 (
            .O(N__40857),
            .I(N__40852));
    LocalMux I__8831 (
            .O(N__40852),
            .I(N__40849));
    Span4Mux_v I__8830 (
            .O(N__40849),
            .I(N__40845));
    InMux I__8829 (
            .O(N__40848),
            .I(N__40842));
    Span4Mux_v I__8828 (
            .O(N__40845),
            .I(N__40839));
    LocalMux I__8827 (
            .O(N__40842),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8826 (
            .O(N__40839),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8825 (
            .O(N__40834),
            .I(N__40828));
    InMux I__8824 (
            .O(N__40833),
            .I(N__40828));
    LocalMux I__8823 (
            .O(N__40828),
            .I(N__40824));
    InMux I__8822 (
            .O(N__40827),
            .I(N__40821));
    Span4Mux_v I__8821 (
            .O(N__40824),
            .I(N__40818));
    LocalMux I__8820 (
            .O(N__40821),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__8819 (
            .O(N__40818),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8818 (
            .O(N__40813),
            .I(N__40810));
    LocalMux I__8817 (
            .O(N__40810),
            .I(N__40807));
    Odrv4 I__8816 (
            .O(N__40807),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__8815 (
            .O(N__40804),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__8814 (
            .O(N__40801),
            .I(N__40795));
    InMux I__8813 (
            .O(N__40800),
            .I(N__40795));
    LocalMux I__8812 (
            .O(N__40795),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__8811 (
            .O(N__40792),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__8810 (
            .O(N__40789),
            .I(N__40783));
    InMux I__8809 (
            .O(N__40788),
            .I(N__40779));
    InMux I__8808 (
            .O(N__40787),
            .I(N__40774));
    InMux I__8807 (
            .O(N__40786),
            .I(N__40774));
    LocalMux I__8806 (
            .O(N__40783),
            .I(N__40771));
    InMux I__8805 (
            .O(N__40782),
            .I(N__40768));
    LocalMux I__8804 (
            .O(N__40779),
            .I(N__40763));
    LocalMux I__8803 (
            .O(N__40774),
            .I(N__40763));
    Span4Mux_v I__8802 (
            .O(N__40771),
            .I(N__40758));
    LocalMux I__8801 (
            .O(N__40768),
            .I(N__40758));
    Span4Mux_v I__8800 (
            .O(N__40763),
            .I(N__40748));
    Span4Mux_v I__8799 (
            .O(N__40758),
            .I(N__40745));
    CascadeMux I__8798 (
            .O(N__40757),
            .I(N__40741));
    CascadeMux I__8797 (
            .O(N__40756),
            .I(N__40737));
    CascadeMux I__8796 (
            .O(N__40755),
            .I(N__40733));
    CascadeMux I__8795 (
            .O(N__40754),
            .I(N__40729));
    CascadeMux I__8794 (
            .O(N__40753),
            .I(N__40725));
    CascadeMux I__8793 (
            .O(N__40752),
            .I(N__40721));
    CascadeMux I__8792 (
            .O(N__40751),
            .I(N__40717));
    Span4Mux_h I__8791 (
            .O(N__40748),
            .I(N__40707));
    Span4Mux_h I__8790 (
            .O(N__40745),
            .I(N__40707));
    InMux I__8789 (
            .O(N__40744),
            .I(N__40692));
    InMux I__8788 (
            .O(N__40741),
            .I(N__40692));
    InMux I__8787 (
            .O(N__40740),
            .I(N__40692));
    InMux I__8786 (
            .O(N__40737),
            .I(N__40692));
    InMux I__8785 (
            .O(N__40736),
            .I(N__40692));
    InMux I__8784 (
            .O(N__40733),
            .I(N__40692));
    InMux I__8783 (
            .O(N__40732),
            .I(N__40692));
    InMux I__8782 (
            .O(N__40729),
            .I(N__40675));
    InMux I__8781 (
            .O(N__40728),
            .I(N__40675));
    InMux I__8780 (
            .O(N__40725),
            .I(N__40675));
    InMux I__8779 (
            .O(N__40724),
            .I(N__40675));
    InMux I__8778 (
            .O(N__40721),
            .I(N__40675));
    InMux I__8777 (
            .O(N__40720),
            .I(N__40675));
    InMux I__8776 (
            .O(N__40717),
            .I(N__40675));
    InMux I__8775 (
            .O(N__40716),
            .I(N__40675));
    CascadeMux I__8774 (
            .O(N__40715),
            .I(N__40672));
    CascadeMux I__8773 (
            .O(N__40714),
            .I(N__40668));
    CascadeMux I__8772 (
            .O(N__40713),
            .I(N__40664));
    CascadeMux I__8771 (
            .O(N__40712),
            .I(N__40660));
    Span4Mux_h I__8770 (
            .O(N__40707),
            .I(N__40648));
    LocalMux I__8769 (
            .O(N__40692),
            .I(N__40648));
    LocalMux I__8768 (
            .O(N__40675),
            .I(N__40648));
    InMux I__8767 (
            .O(N__40672),
            .I(N__40631));
    InMux I__8766 (
            .O(N__40671),
            .I(N__40631));
    InMux I__8765 (
            .O(N__40668),
            .I(N__40631));
    InMux I__8764 (
            .O(N__40667),
            .I(N__40631));
    InMux I__8763 (
            .O(N__40664),
            .I(N__40631));
    InMux I__8762 (
            .O(N__40663),
            .I(N__40631));
    InMux I__8761 (
            .O(N__40660),
            .I(N__40631));
    InMux I__8760 (
            .O(N__40659),
            .I(N__40631));
    CascadeMux I__8759 (
            .O(N__40658),
            .I(N__40627));
    CascadeMux I__8758 (
            .O(N__40657),
            .I(N__40623));
    CascadeMux I__8757 (
            .O(N__40656),
            .I(N__40619));
    InMux I__8756 (
            .O(N__40655),
            .I(N__40613));
    Span4Mux_v I__8755 (
            .O(N__40648),
            .I(N__40600));
    LocalMux I__8754 (
            .O(N__40631),
            .I(N__40600));
    InMux I__8753 (
            .O(N__40630),
            .I(N__40585));
    InMux I__8752 (
            .O(N__40627),
            .I(N__40585));
    InMux I__8751 (
            .O(N__40626),
            .I(N__40585));
    InMux I__8750 (
            .O(N__40623),
            .I(N__40585));
    InMux I__8749 (
            .O(N__40622),
            .I(N__40585));
    InMux I__8748 (
            .O(N__40619),
            .I(N__40585));
    InMux I__8747 (
            .O(N__40618),
            .I(N__40585));
    InMux I__8746 (
            .O(N__40617),
            .I(N__40580));
    InMux I__8745 (
            .O(N__40616),
            .I(N__40580));
    LocalMux I__8744 (
            .O(N__40613),
            .I(N__40566));
    InMux I__8743 (
            .O(N__40612),
            .I(N__40563));
    InMux I__8742 (
            .O(N__40611),
            .I(N__40556));
    InMux I__8741 (
            .O(N__40610),
            .I(N__40556));
    InMux I__8740 (
            .O(N__40609),
            .I(N__40556));
    InMux I__8739 (
            .O(N__40608),
            .I(N__40547));
    InMux I__8738 (
            .O(N__40607),
            .I(N__40547));
    InMux I__8737 (
            .O(N__40606),
            .I(N__40547));
    InMux I__8736 (
            .O(N__40605),
            .I(N__40547));
    Span4Mux_h I__8735 (
            .O(N__40600),
            .I(N__40539));
    LocalMux I__8734 (
            .O(N__40585),
            .I(N__40539));
    LocalMux I__8733 (
            .O(N__40580),
            .I(N__40539));
    InMux I__8732 (
            .O(N__40579),
            .I(N__40534));
    InMux I__8731 (
            .O(N__40578),
            .I(N__40534));
    InMux I__8730 (
            .O(N__40577),
            .I(N__40531));
    InMux I__8729 (
            .O(N__40576),
            .I(N__40528));
    InMux I__8728 (
            .O(N__40575),
            .I(N__40521));
    InMux I__8727 (
            .O(N__40574),
            .I(N__40521));
    InMux I__8726 (
            .O(N__40573),
            .I(N__40521));
    InMux I__8725 (
            .O(N__40572),
            .I(N__40512));
    InMux I__8724 (
            .O(N__40571),
            .I(N__40512));
    InMux I__8723 (
            .O(N__40570),
            .I(N__40512));
    InMux I__8722 (
            .O(N__40569),
            .I(N__40512));
    Span4Mux_v I__8721 (
            .O(N__40566),
            .I(N__40506));
    LocalMux I__8720 (
            .O(N__40563),
            .I(N__40506));
    LocalMux I__8719 (
            .O(N__40556),
            .I(N__40501));
    LocalMux I__8718 (
            .O(N__40547),
            .I(N__40501));
    InMux I__8717 (
            .O(N__40546),
            .I(N__40498));
    Span4Mux_v I__8716 (
            .O(N__40539),
            .I(N__40494));
    LocalMux I__8715 (
            .O(N__40534),
            .I(N__40489));
    LocalMux I__8714 (
            .O(N__40531),
            .I(N__40489));
    LocalMux I__8713 (
            .O(N__40528),
            .I(N__40482));
    LocalMux I__8712 (
            .O(N__40521),
            .I(N__40482));
    LocalMux I__8711 (
            .O(N__40512),
            .I(N__40482));
    InMux I__8710 (
            .O(N__40511),
            .I(N__40479));
    Span4Mux_v I__8709 (
            .O(N__40506),
            .I(N__40475));
    Span4Mux_v I__8708 (
            .O(N__40501),
            .I(N__40470));
    LocalMux I__8707 (
            .O(N__40498),
            .I(N__40470));
    CascadeMux I__8706 (
            .O(N__40497),
            .I(N__40466));
    Span4Mux_v I__8705 (
            .O(N__40494),
            .I(N__40462));
    Span12Mux_s11_h I__8704 (
            .O(N__40489),
            .I(N__40459));
    Span4Mux_v I__8703 (
            .O(N__40482),
            .I(N__40456));
    LocalMux I__8702 (
            .O(N__40479),
            .I(N__40453));
    InMux I__8701 (
            .O(N__40478),
            .I(N__40450));
    Span4Mux_s0_v I__8700 (
            .O(N__40475),
            .I(N__40445));
    Span4Mux_v I__8699 (
            .O(N__40470),
            .I(N__40445));
    InMux I__8698 (
            .O(N__40469),
            .I(N__40438));
    InMux I__8697 (
            .O(N__40466),
            .I(N__40438));
    InMux I__8696 (
            .O(N__40465),
            .I(N__40438));
    Span4Mux_v I__8695 (
            .O(N__40462),
            .I(N__40435));
    Span12Mux_v I__8694 (
            .O(N__40459),
            .I(N__40432));
    Span4Mux_v I__8693 (
            .O(N__40456),
            .I(N__40427));
    Span4Mux_v I__8692 (
            .O(N__40453),
            .I(N__40427));
    LocalMux I__8691 (
            .O(N__40450),
            .I(N__40422));
    Sp12to4 I__8690 (
            .O(N__40445),
            .I(N__40422));
    LocalMux I__8689 (
            .O(N__40438),
            .I(N__40419));
    Span4Mux_h I__8688 (
            .O(N__40435),
            .I(N__40416));
    Span12Mux_v I__8687 (
            .O(N__40432),
            .I(N__40409));
    Sp12to4 I__8686 (
            .O(N__40427),
            .I(N__40409));
    Span12Mux_s11_h I__8685 (
            .O(N__40422),
            .I(N__40409));
    Span4Mux_v I__8684 (
            .O(N__40419),
            .I(N__40406));
    Odrv4 I__8683 (
            .O(N__40416),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__8682 (
            .O(N__40409),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8681 (
            .O(N__40406),
            .I(CONSTANT_ONE_NET));
    InMux I__8680 (
            .O(N__40399),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__8679 (
            .O(N__40396),
            .I(N__40393));
    LocalMux I__8678 (
            .O(N__40393),
            .I(N__40390));
    Odrv4 I__8677 (
            .O(N__40390),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__8676 (
            .O(N__40387),
            .I(bfn_15_27_0_));
    InMux I__8675 (
            .O(N__40384),
            .I(N__40379));
    InMux I__8674 (
            .O(N__40383),
            .I(N__40376));
    InMux I__8673 (
            .O(N__40382),
            .I(N__40373));
    LocalMux I__8672 (
            .O(N__40379),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__8671 (
            .O(N__40376),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__8670 (
            .O(N__40373),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    CascadeMux I__8669 (
            .O(N__40366),
            .I(N__40362));
    InMux I__8668 (
            .O(N__40365),
            .I(N__40359));
    InMux I__8667 (
            .O(N__40362),
            .I(N__40356));
    LocalMux I__8666 (
            .O(N__40359),
            .I(N__40349));
    LocalMux I__8665 (
            .O(N__40356),
            .I(N__40349));
    InMux I__8664 (
            .O(N__40355),
            .I(N__40346));
    InMux I__8663 (
            .O(N__40354),
            .I(N__40343));
    Span4Mux_v I__8662 (
            .O(N__40349),
            .I(N__40340));
    LocalMux I__8661 (
            .O(N__40346),
            .I(N__40337));
    LocalMux I__8660 (
            .O(N__40343),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__8659 (
            .O(N__40340),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__8658 (
            .O(N__40337),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__8657 (
            .O(N__40330),
            .I(N__40327));
    LocalMux I__8656 (
            .O(N__40327),
            .I(N__40324));
    Span4Mux_v I__8655 (
            .O(N__40324),
            .I(N__40321));
    Span4Mux_h I__8654 (
            .O(N__40321),
            .I(N__40318));
    Sp12to4 I__8653 (
            .O(N__40318),
            .I(N__40314));
    InMux I__8652 (
            .O(N__40317),
            .I(N__40311));
    Odrv12 I__8651 (
            .O(N__40314),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    LocalMux I__8650 (
            .O(N__40311),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__8649 (
            .O(N__40306),
            .I(N__40303));
    LocalMux I__8648 (
            .O(N__40303),
            .I(N__40300));
    Span4Mux_v I__8647 (
            .O(N__40300),
            .I(N__40297));
    Sp12to4 I__8646 (
            .O(N__40297),
            .I(N__40294));
    Span12Mux_h I__8645 (
            .O(N__40294),
            .I(N__40291));
    Odrv12 I__8644 (
            .O(N__40291),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__8643 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__8642 (
            .O(N__40285),
            .I(N__40282));
    Span4Mux_v I__8641 (
            .O(N__40282),
            .I(N__40279));
    Sp12to4 I__8640 (
            .O(N__40279),
            .I(N__40276));
    Odrv12 I__8639 (
            .O(N__40276),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__8638 (
            .O(N__40273),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__8637 (
            .O(N__40270),
            .I(N__40267));
    LocalMux I__8636 (
            .O(N__40267),
            .I(N__40264));
    Sp12to4 I__8635 (
            .O(N__40264),
            .I(N__40261));
    Span12Mux_s6_v I__8634 (
            .O(N__40261),
            .I(N__40258));
    Odrv12 I__8633 (
            .O(N__40258),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__8632 (
            .O(N__40255),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__8631 (
            .O(N__40252),
            .I(N__40249));
    LocalMux I__8630 (
            .O(N__40249),
            .I(N__40246));
    Span12Mux_s6_v I__8629 (
            .O(N__40246),
            .I(N__40243));
    Odrv12 I__8628 (
            .O(N__40243),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__8627 (
            .O(N__40240),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__8626 (
            .O(N__40237),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__8625 (
            .O(N__40234),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    CascadeMux I__8624 (
            .O(N__40231),
            .I(N__40228));
    InMux I__8623 (
            .O(N__40228),
            .I(N__40224));
    InMux I__8622 (
            .O(N__40227),
            .I(N__40221));
    LocalMux I__8621 (
            .O(N__40224),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__8620 (
            .O(N__40221),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__8619 (
            .O(N__40216),
            .I(N__40213));
    LocalMux I__8618 (
            .O(N__40213),
            .I(N__40209));
    InMux I__8617 (
            .O(N__40212),
            .I(N__40206));
    Odrv4 I__8616 (
            .O(N__40209),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__8615 (
            .O(N__40206),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    CascadeMux I__8614 (
            .O(N__40201),
            .I(N__40197));
    InMux I__8613 (
            .O(N__40200),
            .I(N__40194));
    InMux I__8612 (
            .O(N__40197),
            .I(N__40191));
    LocalMux I__8611 (
            .O(N__40194),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__8610 (
            .O(N__40191),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__8609 (
            .O(N__40186),
            .I(N__40183));
    LocalMux I__8608 (
            .O(N__40183),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__8607 (
            .O(N__40180),
            .I(N__40174));
    InMux I__8606 (
            .O(N__40179),
            .I(N__40174));
    LocalMux I__8605 (
            .O(N__40174),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__8604 (
            .O(N__40171),
            .I(N__40168));
    LocalMux I__8603 (
            .O(N__40168),
            .I(N__40164));
    InMux I__8602 (
            .O(N__40167),
            .I(N__40161));
    Odrv4 I__8601 (
            .O(N__40164),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__8600 (
            .O(N__40161),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    CascadeMux I__8599 (
            .O(N__40156),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__8598 (
            .O(N__40153),
            .I(N__40150));
    LocalMux I__8597 (
            .O(N__40150),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__8596 (
            .O(N__40147),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    InMux I__8595 (
            .O(N__40144),
            .I(N__40141));
    LocalMux I__8594 (
            .O(N__40141),
            .I(N__40138));
    Odrv4 I__8593 (
            .O(N__40138),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__8592 (
            .O(N__40135),
            .I(N__40132));
    InMux I__8591 (
            .O(N__40132),
            .I(N__40126));
    InMux I__8590 (
            .O(N__40131),
            .I(N__40126));
    LocalMux I__8589 (
            .O(N__40126),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__8588 (
            .O(N__40123),
            .I(N__40120));
    LocalMux I__8587 (
            .O(N__40120),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__8586 (
            .O(N__40117),
            .I(N__40114));
    LocalMux I__8585 (
            .O(N__40114),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    CascadeMux I__8584 (
            .O(N__40111),
            .I(N__40108));
    InMux I__8583 (
            .O(N__40108),
            .I(N__40102));
    InMux I__8582 (
            .O(N__40107),
            .I(N__40102));
    LocalMux I__8581 (
            .O(N__40102),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    CascadeMux I__8580 (
            .O(N__40099),
            .I(N__40095));
    InMux I__8579 (
            .O(N__40098),
            .I(N__40090));
    InMux I__8578 (
            .O(N__40095),
            .I(N__40090));
    LocalMux I__8577 (
            .O(N__40090),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__8576 (
            .O(N__40087),
            .I(N__40084));
    LocalMux I__8575 (
            .O(N__40084),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__8574 (
            .O(N__40081),
            .I(N__40075));
    InMux I__8573 (
            .O(N__40080),
            .I(N__40075));
    LocalMux I__8572 (
            .O(N__40075),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__8571 (
            .O(N__40072),
            .I(N__40068));
    InMux I__8570 (
            .O(N__40071),
            .I(N__40065));
    LocalMux I__8569 (
            .O(N__40068),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__8568 (
            .O(N__40065),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    CascadeMux I__8567 (
            .O(N__40060),
            .I(N__40057));
    InMux I__8566 (
            .O(N__40057),
            .I(N__40051));
    InMux I__8565 (
            .O(N__40056),
            .I(N__40051));
    LocalMux I__8564 (
            .O(N__40051),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__8563 (
            .O(N__40048),
            .I(N__40044));
    InMux I__8562 (
            .O(N__40047),
            .I(N__40041));
    LocalMux I__8561 (
            .O(N__40044),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__8560 (
            .O(N__40041),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    CascadeMux I__8559 (
            .O(N__40036),
            .I(N__40032));
    InMux I__8558 (
            .O(N__40035),
            .I(N__40028));
    InMux I__8557 (
            .O(N__40032),
            .I(N__40023));
    InMux I__8556 (
            .O(N__40031),
            .I(N__40023));
    LocalMux I__8555 (
            .O(N__40028),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__8554 (
            .O(N__40023),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__8553 (
            .O(N__40018),
            .I(N__40015));
    InMux I__8552 (
            .O(N__40015),
            .I(N__40010));
    InMux I__8551 (
            .O(N__40014),
            .I(N__40005));
    InMux I__8550 (
            .O(N__40013),
            .I(N__40005));
    LocalMux I__8549 (
            .O(N__40010),
            .I(N__40000));
    LocalMux I__8548 (
            .O(N__40005),
            .I(N__40000));
    Span4Mux_h I__8547 (
            .O(N__40000),
            .I(N__39997));
    Span4Mux_v I__8546 (
            .O(N__39997),
            .I(N__39993));
    InMux I__8545 (
            .O(N__39996),
            .I(N__39990));
    Span4Mux_v I__8544 (
            .O(N__39993),
            .I(N__39987));
    LocalMux I__8543 (
            .O(N__39990),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__8542 (
            .O(N__39987),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__8541 (
            .O(N__39982),
            .I(N__39978));
    InMux I__8540 (
            .O(N__39981),
            .I(N__39975));
    LocalMux I__8539 (
            .O(N__39978),
            .I(N__39972));
    LocalMux I__8538 (
            .O(N__39975),
            .I(N__39969));
    Span4Mux_h I__8537 (
            .O(N__39972),
            .I(N__39966));
    Span4Mux_s3_h I__8536 (
            .O(N__39969),
            .I(N__39963));
    Span4Mux_h I__8535 (
            .O(N__39966),
            .I(N__39960));
    Span4Mux_h I__8534 (
            .O(N__39963),
            .I(N__39957));
    Odrv4 I__8533 (
            .O(N__39960),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__8532 (
            .O(N__39957),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__8531 (
            .O(N__39952),
            .I(N__39949));
    LocalMux I__8530 (
            .O(N__39949),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__8529 (
            .O(N__39946),
            .I(N__39943));
    InMux I__8528 (
            .O(N__39943),
            .I(N__39939));
    CascadeMux I__8527 (
            .O(N__39942),
            .I(N__39936));
    LocalMux I__8526 (
            .O(N__39939),
            .I(N__39933));
    InMux I__8525 (
            .O(N__39936),
            .I(N__39929));
    Span4Mux_v I__8524 (
            .O(N__39933),
            .I(N__39926));
    InMux I__8523 (
            .O(N__39932),
            .I(N__39923));
    LocalMux I__8522 (
            .O(N__39929),
            .I(N__39920));
    Span4Mux_h I__8521 (
            .O(N__39926),
            .I(N__39917));
    LocalMux I__8520 (
            .O(N__39923),
            .I(N__39912));
    Span4Mux_v I__8519 (
            .O(N__39920),
            .I(N__39907));
    Span4Mux_h I__8518 (
            .O(N__39917),
            .I(N__39907));
    InMux I__8517 (
            .O(N__39916),
            .I(N__39904));
    InMux I__8516 (
            .O(N__39915),
            .I(N__39901));
    Span12Mux_v I__8515 (
            .O(N__39912),
            .I(N__39898));
    Span4Mux_v I__8514 (
            .O(N__39907),
            .I(N__39893));
    LocalMux I__8513 (
            .O(N__39904),
            .I(N__39893));
    LocalMux I__8512 (
            .O(N__39901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__8511 (
            .O(N__39898),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__8510 (
            .O(N__39893),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__8509 (
            .O(N__39886),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__8508 (
            .O(N__39883),
            .I(N__39877));
    InMux I__8507 (
            .O(N__39882),
            .I(N__39877));
    LocalMux I__8506 (
            .O(N__39877),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__8505 (
            .O(N__39874),
            .I(N__39868));
    InMux I__8504 (
            .O(N__39873),
            .I(N__39868));
    LocalMux I__8503 (
            .O(N__39868),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__8502 (
            .O(N__39865),
            .I(N__39859));
    InMux I__8501 (
            .O(N__39864),
            .I(N__39859));
    LocalMux I__8500 (
            .O(N__39859),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    CascadeMux I__8499 (
            .O(N__39856),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__8498 (
            .O(N__39853),
            .I(N__39847));
    InMux I__8497 (
            .O(N__39852),
            .I(N__39847));
    LocalMux I__8496 (
            .O(N__39847),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    CascadeMux I__8495 (
            .O(N__39844),
            .I(N__39841));
    InMux I__8494 (
            .O(N__39841),
            .I(N__39837));
    InMux I__8493 (
            .O(N__39840),
            .I(N__39834));
    LocalMux I__8492 (
            .O(N__39837),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__8491 (
            .O(N__39834),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__8490 (
            .O(N__39829),
            .I(N__39823));
    InMux I__8489 (
            .O(N__39828),
            .I(N__39823));
    LocalMux I__8488 (
            .O(N__39823),
            .I(N__39819));
    InMux I__8487 (
            .O(N__39822),
            .I(N__39816));
    Span4Mux_h I__8486 (
            .O(N__39819),
            .I(N__39813));
    LocalMux I__8485 (
            .O(N__39816),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__8484 (
            .O(N__39813),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__8483 (
            .O(N__39808),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    CascadeMux I__8482 (
            .O(N__39805),
            .I(N__39801));
    CascadeMux I__8481 (
            .O(N__39804),
            .I(N__39798));
    InMux I__8480 (
            .O(N__39801),
            .I(N__39793));
    InMux I__8479 (
            .O(N__39798),
            .I(N__39793));
    LocalMux I__8478 (
            .O(N__39793),
            .I(N__39789));
    InMux I__8477 (
            .O(N__39792),
            .I(N__39786));
    Span4Mux_h I__8476 (
            .O(N__39789),
            .I(N__39783));
    LocalMux I__8475 (
            .O(N__39786),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__8474 (
            .O(N__39783),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__8473 (
            .O(N__39778),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__8472 (
            .O(N__39775),
            .I(N__39772));
    InMux I__8471 (
            .O(N__39772),
            .I(N__39766));
    InMux I__8470 (
            .O(N__39771),
            .I(N__39766));
    LocalMux I__8469 (
            .O(N__39766),
            .I(N__39762));
    InMux I__8468 (
            .O(N__39765),
            .I(N__39759));
    Span4Mux_h I__8467 (
            .O(N__39762),
            .I(N__39756));
    LocalMux I__8466 (
            .O(N__39759),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__8465 (
            .O(N__39756),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__8464 (
            .O(N__39751),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__8463 (
            .O(N__39748),
            .I(N__39742));
    InMux I__8462 (
            .O(N__39747),
            .I(N__39742));
    LocalMux I__8461 (
            .O(N__39742),
            .I(N__39738));
    InMux I__8460 (
            .O(N__39741),
            .I(N__39735));
    Span4Mux_h I__8459 (
            .O(N__39738),
            .I(N__39732));
    LocalMux I__8458 (
            .O(N__39735),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__8457 (
            .O(N__39732),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__8456 (
            .O(N__39727),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__8455 (
            .O(N__39724),
            .I(N__39720));
    InMux I__8454 (
            .O(N__39723),
            .I(N__39717));
    InMux I__8453 (
            .O(N__39720),
            .I(N__39714));
    LocalMux I__8452 (
            .O(N__39717),
            .I(N__39708));
    LocalMux I__8451 (
            .O(N__39714),
            .I(N__39708));
    InMux I__8450 (
            .O(N__39713),
            .I(N__39705));
    Span4Mux_h I__8449 (
            .O(N__39708),
            .I(N__39702));
    LocalMux I__8448 (
            .O(N__39705),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__8447 (
            .O(N__39702),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__8446 (
            .O(N__39697),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__8445 (
            .O(N__39694),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__8444 (
            .O(N__39691),
            .I(N__39688));
    InMux I__8443 (
            .O(N__39688),
            .I(N__39684));
    InMux I__8442 (
            .O(N__39687),
            .I(N__39681));
    LocalMux I__8441 (
            .O(N__39684),
            .I(N__39677));
    LocalMux I__8440 (
            .O(N__39681),
            .I(N__39674));
    InMux I__8439 (
            .O(N__39680),
            .I(N__39671));
    Span4Mux_v I__8438 (
            .O(N__39677),
            .I(N__39668));
    Span12Mux_v I__8437 (
            .O(N__39674),
            .I(N__39665));
    LocalMux I__8436 (
            .O(N__39671),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__8435 (
            .O(N__39668),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__8434 (
            .O(N__39665),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__8433 (
            .O(N__39658),
            .I(N__39655));
    LocalMux I__8432 (
            .O(N__39655),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__8431 (
            .O(N__39652),
            .I(bfn_15_14_0_));
    InMux I__8430 (
            .O(N__39649),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__8429 (
            .O(N__39646),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__8428 (
            .O(N__39643),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__8427 (
            .O(N__39640),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__8426 (
            .O(N__39637),
            .I(N__39631));
    InMux I__8425 (
            .O(N__39636),
            .I(N__39631));
    LocalMux I__8424 (
            .O(N__39631),
            .I(N__39627));
    InMux I__8423 (
            .O(N__39630),
            .I(N__39624));
    Span4Mux_v I__8422 (
            .O(N__39627),
            .I(N__39621));
    LocalMux I__8421 (
            .O(N__39624),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__8420 (
            .O(N__39621),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__8419 (
            .O(N__39616),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    CascadeMux I__8418 (
            .O(N__39613),
            .I(N__39609));
    InMux I__8417 (
            .O(N__39612),
            .I(N__39604));
    InMux I__8416 (
            .O(N__39609),
            .I(N__39604));
    LocalMux I__8415 (
            .O(N__39604),
            .I(N__39600));
    InMux I__8414 (
            .O(N__39603),
            .I(N__39597));
    Span12Mux_s7_v I__8413 (
            .O(N__39600),
            .I(N__39594));
    LocalMux I__8412 (
            .O(N__39597),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv12 I__8411 (
            .O(N__39594),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__8410 (
            .O(N__39589),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__8409 (
            .O(N__39586),
            .I(N__39581));
    InMux I__8408 (
            .O(N__39585),
            .I(N__39576));
    InMux I__8407 (
            .O(N__39584),
            .I(N__39576));
    LocalMux I__8406 (
            .O(N__39581),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__8405 (
            .O(N__39576),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__8404 (
            .O(N__39571),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__8403 (
            .O(N__39568),
            .I(N__39561));
    InMux I__8402 (
            .O(N__39567),
            .I(N__39561));
    InMux I__8401 (
            .O(N__39566),
            .I(N__39558));
    LocalMux I__8400 (
            .O(N__39561),
            .I(N__39555));
    LocalMux I__8399 (
            .O(N__39558),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__8398 (
            .O(N__39555),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__8397 (
            .O(N__39550),
            .I(bfn_15_15_0_));
    InMux I__8396 (
            .O(N__39547),
            .I(N__39543));
    InMux I__8395 (
            .O(N__39546),
            .I(N__39540));
    LocalMux I__8394 (
            .O(N__39543),
            .I(N__39537));
    LocalMux I__8393 (
            .O(N__39540),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__8392 (
            .O(N__39537),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8391 (
            .O(N__39532),
            .I(bfn_15_13_0_));
    InMux I__8390 (
            .O(N__39529),
            .I(N__39525));
    InMux I__8389 (
            .O(N__39528),
            .I(N__39522));
    LocalMux I__8388 (
            .O(N__39525),
            .I(N__39519));
    LocalMux I__8387 (
            .O(N__39522),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__8386 (
            .O(N__39519),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8385 (
            .O(N__39514),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__8384 (
            .O(N__39511),
            .I(N__39507));
    InMux I__8383 (
            .O(N__39510),
            .I(N__39504));
    LocalMux I__8382 (
            .O(N__39507),
            .I(N__39501));
    LocalMux I__8381 (
            .O(N__39504),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__8380 (
            .O(N__39501),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8379 (
            .O(N__39496),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__8378 (
            .O(N__39493),
            .I(N__39489));
    InMux I__8377 (
            .O(N__39492),
            .I(N__39486));
    LocalMux I__8376 (
            .O(N__39489),
            .I(N__39483));
    LocalMux I__8375 (
            .O(N__39486),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__8374 (
            .O(N__39483),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8373 (
            .O(N__39478),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__8372 (
            .O(N__39475),
            .I(N__39471));
    InMux I__8371 (
            .O(N__39474),
            .I(N__39468));
    LocalMux I__8370 (
            .O(N__39471),
            .I(N__39465));
    LocalMux I__8369 (
            .O(N__39468),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__8368 (
            .O(N__39465),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8367 (
            .O(N__39460),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__8366 (
            .O(N__39457),
            .I(N__39454));
    LocalMux I__8365 (
            .O(N__39454),
            .I(N__39450));
    InMux I__8364 (
            .O(N__39453),
            .I(N__39447));
    Span4Mux_v I__8363 (
            .O(N__39450),
            .I(N__39444));
    LocalMux I__8362 (
            .O(N__39447),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__8361 (
            .O(N__39444),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8360 (
            .O(N__39439),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__8359 (
            .O(N__39436),
            .I(N__39432));
    InMux I__8358 (
            .O(N__39435),
            .I(N__39429));
    LocalMux I__8357 (
            .O(N__39432),
            .I(N__39426));
    LocalMux I__8356 (
            .O(N__39429),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__8355 (
            .O(N__39426),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8354 (
            .O(N__39421),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__8353 (
            .O(N__39418),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__8352 (
            .O(N__39415),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__8351 (
            .O(N__39412),
            .I(N__39409));
    InMux I__8350 (
            .O(N__39409),
            .I(N__39404));
    InMux I__8349 (
            .O(N__39408),
            .I(N__39401));
    CascadeMux I__8348 (
            .O(N__39407),
            .I(N__39398));
    LocalMux I__8347 (
            .O(N__39404),
            .I(N__39393));
    LocalMux I__8346 (
            .O(N__39401),
            .I(N__39393));
    InMux I__8345 (
            .O(N__39398),
            .I(N__39390));
    Span4Mux_v I__8344 (
            .O(N__39393),
            .I(N__39387));
    LocalMux I__8343 (
            .O(N__39390),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8342 (
            .O(N__39387),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8341 (
            .O(N__39382),
            .I(N__39378));
    InMux I__8340 (
            .O(N__39381),
            .I(N__39375));
    LocalMux I__8339 (
            .O(N__39378),
            .I(N__39372));
    LocalMux I__8338 (
            .O(N__39375),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv12 I__8337 (
            .O(N__39372),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8336 (
            .O(N__39367),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__8335 (
            .O(N__39364),
            .I(N__39360));
    InMux I__8334 (
            .O(N__39363),
            .I(N__39357));
    LocalMux I__8333 (
            .O(N__39360),
            .I(N__39354));
    LocalMux I__8332 (
            .O(N__39357),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__8331 (
            .O(N__39354),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8330 (
            .O(N__39349),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__8329 (
            .O(N__39346),
            .I(N__39342));
    InMux I__8328 (
            .O(N__39345),
            .I(N__39339));
    LocalMux I__8327 (
            .O(N__39342),
            .I(N__39336));
    LocalMux I__8326 (
            .O(N__39339),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__8325 (
            .O(N__39336),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8324 (
            .O(N__39331),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__8323 (
            .O(N__39328),
            .I(N__39324));
    InMux I__8322 (
            .O(N__39327),
            .I(N__39321));
    LocalMux I__8321 (
            .O(N__39324),
            .I(N__39318));
    LocalMux I__8320 (
            .O(N__39321),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__8319 (
            .O(N__39318),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8318 (
            .O(N__39313),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__8317 (
            .O(N__39310),
            .I(N__39306));
    InMux I__8316 (
            .O(N__39309),
            .I(N__39303));
    LocalMux I__8315 (
            .O(N__39306),
            .I(N__39300));
    LocalMux I__8314 (
            .O(N__39303),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__8313 (
            .O(N__39300),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8312 (
            .O(N__39295),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__8311 (
            .O(N__39292),
            .I(N__39288));
    InMux I__8310 (
            .O(N__39291),
            .I(N__39285));
    LocalMux I__8309 (
            .O(N__39288),
            .I(N__39282));
    LocalMux I__8308 (
            .O(N__39285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__8307 (
            .O(N__39282),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8306 (
            .O(N__39277),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__8305 (
            .O(N__39274),
            .I(N__39270));
    InMux I__8304 (
            .O(N__39273),
            .I(N__39267));
    LocalMux I__8303 (
            .O(N__39270),
            .I(N__39264));
    LocalMux I__8302 (
            .O(N__39267),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__8301 (
            .O(N__39264),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8300 (
            .O(N__39259),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__8299 (
            .O(N__39256),
            .I(N__39253));
    LocalMux I__8298 (
            .O(N__39253),
            .I(N__39250));
    Odrv12 I__8297 (
            .O(N__39250),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__8296 (
            .O(N__39247),
            .I(N__39244));
    InMux I__8295 (
            .O(N__39244),
            .I(N__39241));
    LocalMux I__8294 (
            .O(N__39241),
            .I(N__39238));
    Span4Mux_v I__8293 (
            .O(N__39238),
            .I(N__39235));
    Odrv4 I__8292 (
            .O(N__39235),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__8291 (
            .O(N__39232),
            .I(N__39229));
    LocalMux I__8290 (
            .O(N__39229),
            .I(N__39226));
    Odrv4 I__8289 (
            .O(N__39226),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    CascadeMux I__8288 (
            .O(N__39223),
            .I(N__39220));
    InMux I__8287 (
            .O(N__39220),
            .I(N__39217));
    LocalMux I__8286 (
            .O(N__39217),
            .I(N__39214));
    Odrv4 I__8285 (
            .O(N__39214),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    InMux I__8284 (
            .O(N__39211),
            .I(N__39208));
    LocalMux I__8283 (
            .O(N__39208),
            .I(N__39205));
    Odrv12 I__8282 (
            .O(N__39205),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__8281 (
            .O(N__39202),
            .I(N__39199));
    InMux I__8280 (
            .O(N__39199),
            .I(N__39196));
    LocalMux I__8279 (
            .O(N__39196),
            .I(N__39193));
    Odrv12 I__8278 (
            .O(N__39193),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__8277 (
            .O(N__39190),
            .I(N__39187));
    LocalMux I__8276 (
            .O(N__39187),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    CascadeMux I__8275 (
            .O(N__39184),
            .I(N__39181));
    InMux I__8274 (
            .O(N__39181),
            .I(N__39178));
    LocalMux I__8273 (
            .O(N__39178),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__8272 (
            .O(N__39175),
            .I(N__39172));
    LocalMux I__8271 (
            .O(N__39172),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    CascadeMux I__8270 (
            .O(N__39169),
            .I(N__39166));
    InMux I__8269 (
            .O(N__39166),
            .I(N__39163));
    LocalMux I__8268 (
            .O(N__39163),
            .I(N__39160));
    Odrv4 I__8267 (
            .O(N__39160),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__8266 (
            .O(N__39157),
            .I(N__39154));
    LocalMux I__8265 (
            .O(N__39154),
            .I(N__39151));
    Span4Mux_v I__8264 (
            .O(N__39151),
            .I(N__39148));
    Odrv4 I__8263 (
            .O(N__39148),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__8262 (
            .O(N__39145),
            .I(N__39142));
    InMux I__8261 (
            .O(N__39142),
            .I(N__39139));
    LocalMux I__8260 (
            .O(N__39139),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__8259 (
            .O(N__39136),
            .I(N__39133));
    LocalMux I__8258 (
            .O(N__39133),
            .I(N__39130));
    Odrv12 I__8257 (
            .O(N__39130),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__8256 (
            .O(N__39127),
            .I(N__39124));
    InMux I__8255 (
            .O(N__39124),
            .I(N__39121));
    LocalMux I__8254 (
            .O(N__39121),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__8253 (
            .O(N__39118),
            .I(N__39115));
    InMux I__8252 (
            .O(N__39115),
            .I(N__39112));
    LocalMux I__8251 (
            .O(N__39112),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__8250 (
            .O(N__39109),
            .I(N__39106));
    InMux I__8249 (
            .O(N__39106),
            .I(N__39103));
    LocalMux I__8248 (
            .O(N__39103),
            .I(N__39100));
    Odrv12 I__8247 (
            .O(N__39100),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8246 (
            .O(N__39097),
            .I(N__39094));
    LocalMux I__8245 (
            .O(N__39094),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8244 (
            .O(N__39091),
            .I(N__39088));
    LocalMux I__8243 (
            .O(N__39088),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__8242 (
            .O(N__39085),
            .I(N__39082));
    InMux I__8241 (
            .O(N__39082),
            .I(N__39079));
    LocalMux I__8240 (
            .O(N__39079),
            .I(N__39076));
    Odrv4 I__8239 (
            .O(N__39076),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__8238 (
            .O(N__39073),
            .I(N__39070));
    LocalMux I__8237 (
            .O(N__39070),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8236 (
            .O(N__39067),
            .I(N__39064));
    InMux I__8235 (
            .O(N__39064),
            .I(N__39061));
    LocalMux I__8234 (
            .O(N__39061),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__8233 (
            .O(N__39058),
            .I(N__39055));
    LocalMux I__8232 (
            .O(N__39055),
            .I(N__39052));
    Odrv12 I__8231 (
            .O(N__39052),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__8230 (
            .O(N__39049),
            .I(N__39046));
    InMux I__8229 (
            .O(N__39046),
            .I(N__39043));
    LocalMux I__8228 (
            .O(N__39043),
            .I(N__39040));
    Odrv4 I__8227 (
            .O(N__39040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__8226 (
            .O(N__39037),
            .I(N__39034));
    LocalMux I__8225 (
            .O(N__39034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__8224 (
            .O(N__39031),
            .I(N__39028));
    InMux I__8223 (
            .O(N__39028),
            .I(N__39025));
    LocalMux I__8222 (
            .O(N__39025),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8221 (
            .O(N__39022),
            .I(N__39019));
    InMux I__8220 (
            .O(N__39019),
            .I(N__39016));
    LocalMux I__8219 (
            .O(N__39016),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__8218 (
            .O(N__39013),
            .I(N__39010));
    LocalMux I__8217 (
            .O(N__39010),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__8216 (
            .O(N__39007),
            .I(N__39004));
    LocalMux I__8215 (
            .O(N__39004),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__8214 (
            .O(N__39001),
            .I(N__38998));
    InMux I__8213 (
            .O(N__38998),
            .I(N__38995));
    LocalMux I__8212 (
            .O(N__38995),
            .I(N__38992));
    Odrv4 I__8211 (
            .O(N__38992),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__8210 (
            .O(N__38989),
            .I(N__38986));
    LocalMux I__8209 (
            .O(N__38986),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__8208 (
            .O(N__38983),
            .I(N__38980));
    InMux I__8207 (
            .O(N__38980),
            .I(N__38977));
    LocalMux I__8206 (
            .O(N__38977),
            .I(N__38974));
    Odrv4 I__8205 (
            .O(N__38974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__8204 (
            .O(N__38971),
            .I(N__38968));
    LocalMux I__8203 (
            .O(N__38968),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__8202 (
            .O(N__38965),
            .I(N__38962));
    InMux I__8201 (
            .O(N__38962),
            .I(N__38959));
    LocalMux I__8200 (
            .O(N__38959),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__8199 (
            .O(N__38956),
            .I(N__38953));
    LocalMux I__8198 (
            .O(N__38953),
            .I(N__38950));
    Odrv12 I__8197 (
            .O(N__38950),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__8196 (
            .O(N__38947),
            .I(N__38944));
    InMux I__8195 (
            .O(N__38944),
            .I(N__38941));
    LocalMux I__8194 (
            .O(N__38941),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__8193 (
            .O(N__38938),
            .I(N__38932));
    InMux I__8192 (
            .O(N__38937),
            .I(N__38932));
    LocalMux I__8191 (
            .O(N__38932),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__8190 (
            .O(N__38929),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ));
    InMux I__8189 (
            .O(N__38926),
            .I(N__38923));
    LocalMux I__8188 (
            .O(N__38923),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    IoInMux I__8187 (
            .O(N__38920),
            .I(N__38917));
    LocalMux I__8186 (
            .O(N__38917),
            .I(N__38914));
    Span4Mux_s2_v I__8185 (
            .O(N__38914),
            .I(N__38911));
    Span4Mux_h I__8184 (
            .O(N__38911),
            .I(N__38908));
    Odrv4 I__8183 (
            .O(N__38908),
            .I(s4_phy_c));
    CascadeMux I__8182 (
            .O(N__38905),
            .I(N__38902));
    InMux I__8181 (
            .O(N__38902),
            .I(N__38896));
    InMux I__8180 (
            .O(N__38901),
            .I(N__38896));
    LocalMux I__8179 (
            .O(N__38896),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__8178 (
            .O(N__38893),
            .I(N__38890));
    LocalMux I__8177 (
            .O(N__38890),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__8176 (
            .O(N__38887),
            .I(N__38884));
    LocalMux I__8175 (
            .O(N__38884),
            .I(\pwm_generator_inst.threshold_2 ));
    CascadeMux I__8174 (
            .O(N__38881),
            .I(N__38878));
    InMux I__8173 (
            .O(N__38878),
            .I(N__38875));
    LocalMux I__8172 (
            .O(N__38875),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    CascadeMux I__8171 (
            .O(N__38872),
            .I(N__38869));
    InMux I__8170 (
            .O(N__38869),
            .I(N__38866));
    LocalMux I__8169 (
            .O(N__38866),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__8168 (
            .O(N__38863),
            .I(N__38860));
    LocalMux I__8167 (
            .O(N__38860),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    CascadeMux I__8166 (
            .O(N__38857),
            .I(N__38854));
    InMux I__8165 (
            .O(N__38854),
            .I(N__38851));
    LocalMux I__8164 (
            .O(N__38851),
            .I(N__38848));
    Odrv4 I__8163 (
            .O(N__38848),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__8162 (
            .O(N__38845),
            .I(N__38842));
    LocalMux I__8161 (
            .O(N__38842),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__8160 (
            .O(N__38839),
            .I(N__38836));
    InMux I__8159 (
            .O(N__38836),
            .I(N__38833));
    LocalMux I__8158 (
            .O(N__38833),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__8157 (
            .O(N__38830),
            .I(N__38827));
    LocalMux I__8156 (
            .O(N__38827),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__8155 (
            .O(N__38824),
            .I(N__38821));
    LocalMux I__8154 (
            .O(N__38821),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__8153 (
            .O(N__38818),
            .I(N__38815));
    LocalMux I__8152 (
            .O(N__38815),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__8151 (
            .O(N__38812),
            .I(N__38809));
    LocalMux I__8150 (
            .O(N__38809),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__8149 (
            .O(N__38806),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__8148 (
            .O(N__38803),
            .I(N__38794));
    InMux I__8147 (
            .O(N__38802),
            .I(N__38794));
    InMux I__8146 (
            .O(N__38801),
            .I(N__38787));
    InMux I__8145 (
            .O(N__38800),
            .I(N__38774));
    InMux I__8144 (
            .O(N__38799),
            .I(N__38771));
    LocalMux I__8143 (
            .O(N__38794),
            .I(N__38768));
    InMux I__8142 (
            .O(N__38793),
            .I(N__38759));
    InMux I__8141 (
            .O(N__38792),
            .I(N__38759));
    InMux I__8140 (
            .O(N__38791),
            .I(N__38759));
    InMux I__8139 (
            .O(N__38790),
            .I(N__38759));
    LocalMux I__8138 (
            .O(N__38787),
            .I(N__38756));
    InMux I__8137 (
            .O(N__38786),
            .I(N__38745));
    InMux I__8136 (
            .O(N__38785),
            .I(N__38745));
    InMux I__8135 (
            .O(N__38784),
            .I(N__38745));
    InMux I__8134 (
            .O(N__38783),
            .I(N__38745));
    InMux I__8133 (
            .O(N__38782),
            .I(N__38745));
    InMux I__8132 (
            .O(N__38781),
            .I(N__38742));
    InMux I__8131 (
            .O(N__38780),
            .I(N__38739));
    InMux I__8130 (
            .O(N__38779),
            .I(N__38721));
    InMux I__8129 (
            .O(N__38778),
            .I(N__38721));
    InMux I__8128 (
            .O(N__38777),
            .I(N__38721));
    LocalMux I__8127 (
            .O(N__38774),
            .I(N__38712));
    LocalMux I__8126 (
            .O(N__38771),
            .I(N__38712));
    Span4Mux_h I__8125 (
            .O(N__38768),
            .I(N__38712));
    LocalMux I__8124 (
            .O(N__38759),
            .I(N__38712));
    Sp12to4 I__8123 (
            .O(N__38756),
            .I(N__38709));
    LocalMux I__8122 (
            .O(N__38745),
            .I(N__38703));
    LocalMux I__8121 (
            .O(N__38742),
            .I(N__38703));
    LocalMux I__8120 (
            .O(N__38739),
            .I(N__38700));
    InMux I__8119 (
            .O(N__38738),
            .I(N__38694));
    InMux I__8118 (
            .O(N__38737),
            .I(N__38694));
    InMux I__8117 (
            .O(N__38736),
            .I(N__38683));
    InMux I__8116 (
            .O(N__38735),
            .I(N__38683));
    InMux I__8115 (
            .O(N__38734),
            .I(N__38683));
    InMux I__8114 (
            .O(N__38733),
            .I(N__38683));
    InMux I__8113 (
            .O(N__38732),
            .I(N__38683));
    InMux I__8112 (
            .O(N__38731),
            .I(N__38674));
    InMux I__8111 (
            .O(N__38730),
            .I(N__38674));
    InMux I__8110 (
            .O(N__38729),
            .I(N__38674));
    InMux I__8109 (
            .O(N__38728),
            .I(N__38674));
    LocalMux I__8108 (
            .O(N__38721),
            .I(N__38671));
    Span4Mux_v I__8107 (
            .O(N__38712),
            .I(N__38668));
    Span12Mux_h I__8106 (
            .O(N__38709),
            .I(N__38665));
    InMux I__8105 (
            .O(N__38708),
            .I(N__38662));
    Span4Mux_h I__8104 (
            .O(N__38703),
            .I(N__38657));
    Span4Mux_h I__8103 (
            .O(N__38700),
            .I(N__38657));
    InMux I__8102 (
            .O(N__38699),
            .I(N__38654));
    LocalMux I__8101 (
            .O(N__38694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__8100 (
            .O(N__38683),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__8099 (
            .O(N__38674),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__8098 (
            .O(N__38671),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__8097 (
            .O(N__38668),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__8096 (
            .O(N__38665),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__8095 (
            .O(N__38662),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__8094 (
            .O(N__38657),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__8093 (
            .O(N__38654),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__8092 (
            .O(N__38635),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__8091 (
            .O(N__38632),
            .I(N__38629));
    LocalMux I__8090 (
            .O(N__38629),
            .I(N__38626));
    Span4Mux_h I__8089 (
            .O(N__38626),
            .I(N__38623));
    Span4Mux_h I__8088 (
            .O(N__38623),
            .I(N__38620));
    Odrv4 I__8087 (
            .O(N__38620),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__8086 (
            .O(N__38617),
            .I(N__38614));
    LocalMux I__8085 (
            .O(N__38614),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    CascadeMux I__8084 (
            .O(N__38611),
            .I(N__38608));
    InMux I__8083 (
            .O(N__38608),
            .I(N__38605));
    LocalMux I__8082 (
            .O(N__38605),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    CascadeMux I__8081 (
            .O(N__38602),
            .I(N__38599));
    InMux I__8080 (
            .O(N__38599),
            .I(N__38596));
    LocalMux I__8079 (
            .O(N__38596),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__8078 (
            .O(N__38593),
            .I(N__38590));
    LocalMux I__8077 (
            .O(N__38590),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__8076 (
            .O(N__38587),
            .I(N__38584));
    LocalMux I__8075 (
            .O(N__38584),
            .I(\pwm_generator_inst.threshold_4 ));
    CascadeMux I__8074 (
            .O(N__38581),
            .I(N__38578));
    InMux I__8073 (
            .O(N__38578),
            .I(N__38575));
    LocalMux I__8072 (
            .O(N__38575),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    CascadeMux I__8071 (
            .O(N__38572),
            .I(N__38569));
    InMux I__8070 (
            .O(N__38569),
            .I(N__38566));
    LocalMux I__8069 (
            .O(N__38566),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__8068 (
            .O(N__38563),
            .I(N__38560));
    LocalMux I__8067 (
            .O(N__38560),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__8066 (
            .O(N__38557),
            .I(N__38554));
    LocalMux I__8065 (
            .O(N__38554),
            .I(\pwm_generator_inst.un14_counter_1 ));
    CascadeMux I__8064 (
            .O(N__38551),
            .I(N__38548));
    InMux I__8063 (
            .O(N__38548),
            .I(N__38545));
    LocalMux I__8062 (
            .O(N__38545),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    CascadeMux I__8061 (
            .O(N__38542),
            .I(N__38539));
    InMux I__8060 (
            .O(N__38539),
            .I(N__38536));
    LocalMux I__8059 (
            .O(N__38536),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__8058 (
            .O(N__38533),
            .I(N__38530));
    LocalMux I__8057 (
            .O(N__38530),
            .I(N__38527));
    Span4Mux_v I__8056 (
            .O(N__38527),
            .I(N__38524));
    Odrv4 I__8055 (
            .O(N__38524),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__8054 (
            .O(N__38521),
            .I(N__38518));
    InMux I__8053 (
            .O(N__38518),
            .I(N__38515));
    LocalMux I__8052 (
            .O(N__38515),
            .I(N__38512));
    Span4Mux_v I__8051 (
            .O(N__38512),
            .I(N__38508));
    InMux I__8050 (
            .O(N__38511),
            .I(N__38505));
    Span4Mux_v I__8049 (
            .O(N__38508),
            .I(N__38500));
    LocalMux I__8048 (
            .O(N__38505),
            .I(N__38497));
    InMux I__8047 (
            .O(N__38504),
            .I(N__38494));
    InMux I__8046 (
            .O(N__38503),
            .I(N__38491));
    Sp12to4 I__8045 (
            .O(N__38500),
            .I(N__38488));
    Span4Mux_v I__8044 (
            .O(N__38497),
            .I(N__38485));
    LocalMux I__8043 (
            .O(N__38494),
            .I(N__38482));
    LocalMux I__8042 (
            .O(N__38491),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__8041 (
            .O(N__38488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__8040 (
            .O(N__38485),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__8039 (
            .O(N__38482),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__8038 (
            .O(N__38473),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__8037 (
            .O(N__38470),
            .I(N__38467));
    LocalMux I__8036 (
            .O(N__38467),
            .I(N__38464));
    Odrv4 I__8035 (
            .O(N__38464),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__8034 (
            .O(N__38461),
            .I(N__38458));
    InMux I__8033 (
            .O(N__38458),
            .I(N__38455));
    LocalMux I__8032 (
            .O(N__38455),
            .I(N__38452));
    Span4Mux_h I__8031 (
            .O(N__38452),
            .I(N__38449));
    Span4Mux_h I__8030 (
            .O(N__38449),
            .I(N__38444));
    InMux I__8029 (
            .O(N__38448),
            .I(N__38441));
    CascadeMux I__8028 (
            .O(N__38447),
            .I(N__38438));
    Span4Mux_h I__8027 (
            .O(N__38444),
            .I(N__38434));
    LocalMux I__8026 (
            .O(N__38441),
            .I(N__38431));
    InMux I__8025 (
            .O(N__38438),
            .I(N__38428));
    InMux I__8024 (
            .O(N__38437),
            .I(N__38425));
    Span4Mux_v I__8023 (
            .O(N__38434),
            .I(N__38422));
    Span4Mux_v I__8022 (
            .O(N__38431),
            .I(N__38417));
    LocalMux I__8021 (
            .O(N__38428),
            .I(N__38417));
    LocalMux I__8020 (
            .O(N__38425),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__8019 (
            .O(N__38422),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__8018 (
            .O(N__38417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__8017 (
            .O(N__38410),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__8016 (
            .O(N__38407),
            .I(N__38404));
    LocalMux I__8015 (
            .O(N__38404),
            .I(N__38401));
    Odrv12 I__8014 (
            .O(N__38401),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    CascadeMux I__8013 (
            .O(N__38398),
            .I(N__38395));
    InMux I__8012 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__8011 (
            .O(N__38392),
            .I(N__38389));
    Sp12to4 I__8010 (
            .O(N__38389),
            .I(N__38385));
    InMux I__8009 (
            .O(N__38388),
            .I(N__38380));
    Span12Mux_v I__8008 (
            .O(N__38385),
            .I(N__38377));
    InMux I__8007 (
            .O(N__38384),
            .I(N__38374));
    InMux I__8006 (
            .O(N__38383),
            .I(N__38371));
    LocalMux I__8005 (
            .O(N__38380),
            .I(N__38368));
    Odrv12 I__8004 (
            .O(N__38377),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__8003 (
            .O(N__38374),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__8002 (
            .O(N__38371),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__8001 (
            .O(N__38368),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__8000 (
            .O(N__38359),
            .I(bfn_14_20_0_));
    InMux I__7999 (
            .O(N__38356),
            .I(N__38353));
    LocalMux I__7998 (
            .O(N__38353),
            .I(N__38350));
    Odrv12 I__7997 (
            .O(N__38350),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    CascadeMux I__7996 (
            .O(N__38347),
            .I(N__38344));
    InMux I__7995 (
            .O(N__38344),
            .I(N__38341));
    LocalMux I__7994 (
            .O(N__38341),
            .I(N__38338));
    Span4Mux_v I__7993 (
            .O(N__38338),
            .I(N__38334));
    InMux I__7992 (
            .O(N__38337),
            .I(N__38330));
    Sp12to4 I__7991 (
            .O(N__38334),
            .I(N__38326));
    InMux I__7990 (
            .O(N__38333),
            .I(N__38323));
    LocalMux I__7989 (
            .O(N__38330),
            .I(N__38320));
    InMux I__7988 (
            .O(N__38329),
            .I(N__38317));
    Span12Mux_h I__7987 (
            .O(N__38326),
            .I(N__38314));
    LocalMux I__7986 (
            .O(N__38323),
            .I(N__38311));
    Span4Mux_v I__7985 (
            .O(N__38320),
            .I(N__38308));
    LocalMux I__7984 (
            .O(N__38317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__7983 (
            .O(N__38314),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__7982 (
            .O(N__38311),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__7981 (
            .O(N__38308),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__7980 (
            .O(N__38299),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__7979 (
            .O(N__38296),
            .I(N__38293));
    LocalMux I__7978 (
            .O(N__38293),
            .I(N__38290));
    Span4Mux_h I__7977 (
            .O(N__38290),
            .I(N__38287));
    Span4Mux_h I__7976 (
            .O(N__38287),
            .I(N__38284));
    Odrv4 I__7975 (
            .O(N__38284),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    CascadeMux I__7974 (
            .O(N__38281),
            .I(N__38278));
    InMux I__7973 (
            .O(N__38278),
            .I(N__38275));
    LocalMux I__7972 (
            .O(N__38275),
            .I(N__38272));
    Span4Mux_v I__7971 (
            .O(N__38272),
            .I(N__38268));
    CascadeMux I__7970 (
            .O(N__38271),
            .I(N__38265));
    Span4Mux_h I__7969 (
            .O(N__38268),
            .I(N__38261));
    InMux I__7968 (
            .O(N__38265),
            .I(N__38258));
    CascadeMux I__7967 (
            .O(N__38264),
            .I(N__38254));
    Span4Mux_h I__7966 (
            .O(N__38261),
            .I(N__38249));
    LocalMux I__7965 (
            .O(N__38258),
            .I(N__38249));
    InMux I__7964 (
            .O(N__38257),
            .I(N__38246));
    InMux I__7963 (
            .O(N__38254),
            .I(N__38243));
    Span4Mux_h I__7962 (
            .O(N__38249),
            .I(N__38240));
    LocalMux I__7961 (
            .O(N__38246),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__7960 (
            .O(N__38243),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__7959 (
            .O(N__38240),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__7958 (
            .O(N__38233),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__7957 (
            .O(N__38230),
            .I(N__38227));
    LocalMux I__7956 (
            .O(N__38227),
            .I(N__38224));
    Span4Mux_v I__7955 (
            .O(N__38224),
            .I(N__38221));
    Span4Mux_h I__7954 (
            .O(N__38221),
            .I(N__38217));
    InMux I__7953 (
            .O(N__38220),
            .I(N__38214));
    Span4Mux_h I__7952 (
            .O(N__38217),
            .I(N__38207));
    LocalMux I__7951 (
            .O(N__38214),
            .I(N__38207));
    InMux I__7950 (
            .O(N__38213),
            .I(N__38204));
    InMux I__7949 (
            .O(N__38212),
            .I(N__38201));
    Span4Mux_h I__7948 (
            .O(N__38207),
            .I(N__38198));
    LocalMux I__7947 (
            .O(N__38204),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__7946 (
            .O(N__38201),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__7945 (
            .O(N__38198),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__7944 (
            .O(N__38191),
            .I(N__38188));
    InMux I__7943 (
            .O(N__38188),
            .I(N__38185));
    LocalMux I__7942 (
            .O(N__38185),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    InMux I__7941 (
            .O(N__38182),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__7940 (
            .O(N__38179),
            .I(N__38176));
    LocalMux I__7939 (
            .O(N__38176),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    CascadeMux I__7938 (
            .O(N__38173),
            .I(N__38170));
    InMux I__7937 (
            .O(N__38170),
            .I(N__38167));
    LocalMux I__7936 (
            .O(N__38167),
            .I(N__38164));
    Span4Mux_v I__7935 (
            .O(N__38164),
            .I(N__38161));
    Span4Mux_h I__7934 (
            .O(N__38161),
            .I(N__38158));
    Span4Mux_h I__7933 (
            .O(N__38158),
            .I(N__38153));
    InMux I__7932 (
            .O(N__38157),
            .I(N__38149));
    InMux I__7931 (
            .O(N__38156),
            .I(N__38146));
    Span4Mux_h I__7930 (
            .O(N__38153),
            .I(N__38143));
    InMux I__7929 (
            .O(N__38152),
            .I(N__38140));
    LocalMux I__7928 (
            .O(N__38149),
            .I(N__38137));
    LocalMux I__7927 (
            .O(N__38146),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__7926 (
            .O(N__38143),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__7925 (
            .O(N__38140),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__7924 (
            .O(N__38137),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__7923 (
            .O(N__38128),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__7922 (
            .O(N__38125),
            .I(N__38122));
    LocalMux I__7921 (
            .O(N__38122),
            .I(N__38119));
    Span4Mux_h I__7920 (
            .O(N__38119),
            .I(N__38116));
    Span4Mux_h I__7919 (
            .O(N__38116),
            .I(N__38113));
    Odrv4 I__7918 (
            .O(N__38113),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    CascadeMux I__7917 (
            .O(N__38110),
            .I(N__38107));
    InMux I__7916 (
            .O(N__38107),
            .I(N__38104));
    LocalMux I__7915 (
            .O(N__38104),
            .I(N__38101));
    Span4Mux_v I__7914 (
            .O(N__38101),
            .I(N__38097));
    InMux I__7913 (
            .O(N__38100),
            .I(N__38094));
    Sp12to4 I__7912 (
            .O(N__38097),
            .I(N__38089));
    LocalMux I__7911 (
            .O(N__38094),
            .I(N__38086));
    InMux I__7910 (
            .O(N__38093),
            .I(N__38083));
    InMux I__7909 (
            .O(N__38092),
            .I(N__38080));
    Span12Mux_h I__7908 (
            .O(N__38089),
            .I(N__38077));
    Span4Mux_v I__7907 (
            .O(N__38086),
            .I(N__38074));
    LocalMux I__7906 (
            .O(N__38083),
            .I(N__38071));
    LocalMux I__7905 (
            .O(N__38080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv12 I__7904 (
            .O(N__38077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__7903 (
            .O(N__38074),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__7902 (
            .O(N__38071),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__7901 (
            .O(N__38062),
            .I(N__38059));
    LocalMux I__7900 (
            .O(N__38059),
            .I(N__38056));
    Span4Mux_h I__7899 (
            .O(N__38056),
            .I(N__38053));
    Span4Mux_h I__7898 (
            .O(N__38053),
            .I(N__38050));
    Odrv4 I__7897 (
            .O(N__38050),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__7896 (
            .O(N__38047),
            .I(N__38044));
    InMux I__7895 (
            .O(N__38044),
            .I(N__38041));
    LocalMux I__7894 (
            .O(N__38041),
            .I(N__38037));
    InMux I__7893 (
            .O(N__38040),
            .I(N__38033));
    Span4Mux_h I__7892 (
            .O(N__38037),
            .I(N__38030));
    InMux I__7891 (
            .O(N__38036),
            .I(N__38026));
    LocalMux I__7890 (
            .O(N__38033),
            .I(N__38023));
    Sp12to4 I__7889 (
            .O(N__38030),
            .I(N__38020));
    InMux I__7888 (
            .O(N__38029),
            .I(N__38017));
    LocalMux I__7887 (
            .O(N__38026),
            .I(N__38014));
    Span4Mux_v I__7886 (
            .O(N__38023),
            .I(N__38011));
    Span12Mux_v I__7885 (
            .O(N__38020),
            .I(N__38006));
    LocalMux I__7884 (
            .O(N__38017),
            .I(N__38006));
    Odrv12 I__7883 (
            .O(N__38014),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__7882 (
            .O(N__38011),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv12 I__7881 (
            .O(N__38006),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__7880 (
            .O(N__37999),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__7879 (
            .O(N__37996),
            .I(N__37993));
    LocalMux I__7878 (
            .O(N__37993),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__7877 (
            .O(N__37990),
            .I(N__37987));
    InMux I__7876 (
            .O(N__37987),
            .I(N__37984));
    LocalMux I__7875 (
            .O(N__37984),
            .I(N__37980));
    CascadeMux I__7874 (
            .O(N__37983),
            .I(N__37977));
    Span4Mux_v I__7873 (
            .O(N__37980),
            .I(N__37972));
    InMux I__7872 (
            .O(N__37977),
            .I(N__37969));
    InMux I__7871 (
            .O(N__37976),
            .I(N__37966));
    InMux I__7870 (
            .O(N__37975),
            .I(N__37963));
    Span4Mux_h I__7869 (
            .O(N__37972),
            .I(N__37960));
    LocalMux I__7868 (
            .O(N__37969),
            .I(N__37957));
    LocalMux I__7867 (
            .O(N__37966),
            .I(N__37952));
    LocalMux I__7866 (
            .O(N__37963),
            .I(N__37952));
    Span4Mux_h I__7865 (
            .O(N__37960),
            .I(N__37947));
    Span4Mux_v I__7864 (
            .O(N__37957),
            .I(N__37947));
    Odrv12 I__7863 (
            .O(N__37952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__7862 (
            .O(N__37947),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__7861 (
            .O(N__37942),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__7860 (
            .O(N__37939),
            .I(N__37936));
    LocalMux I__7859 (
            .O(N__37936),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__7858 (
            .O(N__37933),
            .I(N__37930));
    InMux I__7857 (
            .O(N__37930),
            .I(N__37927));
    LocalMux I__7856 (
            .O(N__37927),
            .I(N__37921));
    CascadeMux I__7855 (
            .O(N__37926),
            .I(N__37918));
    InMux I__7854 (
            .O(N__37925),
            .I(N__37915));
    InMux I__7853 (
            .O(N__37924),
            .I(N__37912));
    Span12Mux_v I__7852 (
            .O(N__37921),
            .I(N__37909));
    InMux I__7851 (
            .O(N__37918),
            .I(N__37906));
    LocalMux I__7850 (
            .O(N__37915),
            .I(N__37903));
    LocalMux I__7849 (
            .O(N__37912),
            .I(N__37900));
    Odrv12 I__7848 (
            .O(N__37909),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__7847 (
            .O(N__37906),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv12 I__7846 (
            .O(N__37903),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__7845 (
            .O(N__37900),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__7844 (
            .O(N__37891),
            .I(bfn_14_19_0_));
    InMux I__7843 (
            .O(N__37888),
            .I(N__37885));
    LocalMux I__7842 (
            .O(N__37885),
            .I(N__37882));
    Sp12to4 I__7841 (
            .O(N__37882),
            .I(N__37879));
    Span12Mux_v I__7840 (
            .O(N__37879),
            .I(N__37873));
    InMux I__7839 (
            .O(N__37878),
            .I(N__37870));
    InMux I__7838 (
            .O(N__37877),
            .I(N__37867));
    InMux I__7837 (
            .O(N__37876),
            .I(N__37864));
    Span12Mux_h I__7836 (
            .O(N__37873),
            .I(N__37859));
    LocalMux I__7835 (
            .O(N__37870),
            .I(N__37859));
    LocalMux I__7834 (
            .O(N__37867),
            .I(N__37856));
    LocalMux I__7833 (
            .O(N__37864),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv12 I__7832 (
            .O(N__37859),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__7831 (
            .O(N__37856),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__7830 (
            .O(N__37849),
            .I(N__37846));
    InMux I__7829 (
            .O(N__37846),
            .I(N__37843));
    LocalMux I__7828 (
            .O(N__37843),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__7827 (
            .O(N__37840),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__7826 (
            .O(N__37837),
            .I(N__37834));
    LocalMux I__7825 (
            .O(N__37834),
            .I(N__37831));
    Sp12to4 I__7824 (
            .O(N__37831),
            .I(N__37827));
    InMux I__7823 (
            .O(N__37830),
            .I(N__37824));
    Span12Mux_v I__7822 (
            .O(N__37827),
            .I(N__37819));
    LocalMux I__7821 (
            .O(N__37824),
            .I(N__37816));
    InMux I__7820 (
            .O(N__37823),
            .I(N__37813));
    InMux I__7819 (
            .O(N__37822),
            .I(N__37810));
    Span12Mux_h I__7818 (
            .O(N__37819),
            .I(N__37807));
    Span4Mux_v I__7817 (
            .O(N__37816),
            .I(N__37802));
    LocalMux I__7816 (
            .O(N__37813),
            .I(N__37802));
    LocalMux I__7815 (
            .O(N__37810),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__7814 (
            .O(N__37807),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7813 (
            .O(N__37802),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__7812 (
            .O(N__37795),
            .I(N__37792));
    InMux I__7811 (
            .O(N__37792),
            .I(N__37789));
    LocalMux I__7810 (
            .O(N__37789),
            .I(N__37786));
    Odrv4 I__7809 (
            .O(N__37786),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__7808 (
            .O(N__37783),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__7807 (
            .O(N__37780),
            .I(N__37777));
    LocalMux I__7806 (
            .O(N__37777),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__7805 (
            .O(N__37774),
            .I(N__37771));
    InMux I__7804 (
            .O(N__37771),
            .I(N__37768));
    LocalMux I__7803 (
            .O(N__37768),
            .I(N__37765));
    Span4Mux_v I__7802 (
            .O(N__37765),
            .I(N__37759));
    InMux I__7801 (
            .O(N__37764),
            .I(N__37756));
    InMux I__7800 (
            .O(N__37763),
            .I(N__37753));
    InMux I__7799 (
            .O(N__37762),
            .I(N__37750));
    Sp12to4 I__7798 (
            .O(N__37759),
            .I(N__37747));
    LocalMux I__7797 (
            .O(N__37756),
            .I(N__37742));
    LocalMux I__7796 (
            .O(N__37753),
            .I(N__37742));
    LocalMux I__7795 (
            .O(N__37750),
            .I(N__37739));
    Span12Mux_h I__7794 (
            .O(N__37747),
            .I(N__37736));
    Span4Mux_v I__7793 (
            .O(N__37742),
            .I(N__37733));
    Span4Mux_h I__7792 (
            .O(N__37739),
            .I(N__37730));
    Odrv12 I__7791 (
            .O(N__37736),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__7790 (
            .O(N__37733),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__7789 (
            .O(N__37730),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__7788 (
            .O(N__37723),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__7787 (
            .O(N__37720),
            .I(N__37717));
    LocalMux I__7786 (
            .O(N__37717),
            .I(N__37714));
    Odrv4 I__7785 (
            .O(N__37714),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__7784 (
            .O(N__37711),
            .I(N__37708));
    InMux I__7783 (
            .O(N__37708),
            .I(N__37705));
    LocalMux I__7782 (
            .O(N__37705),
            .I(N__37700));
    InMux I__7781 (
            .O(N__37704),
            .I(N__37696));
    InMux I__7780 (
            .O(N__37703),
            .I(N__37693));
    Span12Mux_v I__7779 (
            .O(N__37700),
            .I(N__37690));
    InMux I__7778 (
            .O(N__37699),
            .I(N__37687));
    LocalMux I__7777 (
            .O(N__37696),
            .I(N__37682));
    LocalMux I__7776 (
            .O(N__37693),
            .I(N__37682));
    Odrv12 I__7775 (
            .O(N__37690),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__7774 (
            .O(N__37687),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__7773 (
            .O(N__37682),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__7772 (
            .O(N__37675),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__7771 (
            .O(N__37672),
            .I(N__37669));
    LocalMux I__7770 (
            .O(N__37669),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__7769 (
            .O(N__37666),
            .I(N__37663));
    InMux I__7768 (
            .O(N__37663),
            .I(N__37660));
    LocalMux I__7767 (
            .O(N__37660),
            .I(N__37657));
    Sp12to4 I__7766 (
            .O(N__37657),
            .I(N__37652));
    CascadeMux I__7765 (
            .O(N__37656),
            .I(N__37649));
    CascadeMux I__7764 (
            .O(N__37655),
            .I(N__37646));
    Span12Mux_v I__7763 (
            .O(N__37652),
            .I(N__37642));
    InMux I__7762 (
            .O(N__37649),
            .I(N__37639));
    InMux I__7761 (
            .O(N__37646),
            .I(N__37636));
    InMux I__7760 (
            .O(N__37645),
            .I(N__37633));
    Span12Mux_h I__7759 (
            .O(N__37642),
            .I(N__37628));
    LocalMux I__7758 (
            .O(N__37639),
            .I(N__37628));
    LocalMux I__7757 (
            .O(N__37636),
            .I(N__37625));
    LocalMux I__7756 (
            .O(N__37633),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__7755 (
            .O(N__37628),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__7754 (
            .O(N__37625),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__7753 (
            .O(N__37618),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__7752 (
            .O(N__37615),
            .I(N__37612));
    LocalMux I__7751 (
            .O(N__37612),
            .I(N__37609));
    Odrv12 I__7750 (
            .O(N__37609),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__7749 (
            .O(N__37606),
            .I(N__37603));
    InMux I__7748 (
            .O(N__37603),
            .I(N__37600));
    LocalMux I__7747 (
            .O(N__37600),
            .I(N__37597));
    Span4Mux_h I__7746 (
            .O(N__37597),
            .I(N__37594));
    Span4Mux_h I__7745 (
            .O(N__37594),
            .I(N__37589));
    InMux I__7744 (
            .O(N__37593),
            .I(N__37586));
    InMux I__7743 (
            .O(N__37592),
            .I(N__37583));
    Span4Mux_v I__7742 (
            .O(N__37589),
            .I(N__37577));
    LocalMux I__7741 (
            .O(N__37586),
            .I(N__37577));
    LocalMux I__7740 (
            .O(N__37583),
            .I(N__37574));
    InMux I__7739 (
            .O(N__37582),
            .I(N__37571));
    Span4Mux_h I__7738 (
            .O(N__37577),
            .I(N__37568));
    Span4Mux_v I__7737 (
            .O(N__37574),
            .I(N__37565));
    LocalMux I__7736 (
            .O(N__37571),
            .I(N__37560));
    Span4Mux_v I__7735 (
            .O(N__37568),
            .I(N__37560));
    Odrv4 I__7734 (
            .O(N__37565),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__7733 (
            .O(N__37560),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__7732 (
            .O(N__37555),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__7731 (
            .O(N__37552),
            .I(N__37549));
    LocalMux I__7730 (
            .O(N__37549),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__7729 (
            .O(N__37546),
            .I(N__37543));
    InMux I__7728 (
            .O(N__37543),
            .I(N__37540));
    LocalMux I__7727 (
            .O(N__37540),
            .I(N__37537));
    Span4Mux_h I__7726 (
            .O(N__37537),
            .I(N__37531));
    InMux I__7725 (
            .O(N__37536),
            .I(N__37528));
    InMux I__7724 (
            .O(N__37535),
            .I(N__37525));
    InMux I__7723 (
            .O(N__37534),
            .I(N__37522));
    Sp12to4 I__7722 (
            .O(N__37531),
            .I(N__37519));
    LocalMux I__7721 (
            .O(N__37528),
            .I(N__37514));
    LocalMux I__7720 (
            .O(N__37525),
            .I(N__37514));
    LocalMux I__7719 (
            .O(N__37522),
            .I(N__37511));
    Span12Mux_v I__7718 (
            .O(N__37519),
            .I(N__37508));
    Span4Mux_v I__7717 (
            .O(N__37514),
            .I(N__37503));
    Span4Mux_h I__7716 (
            .O(N__37511),
            .I(N__37503));
    Odrv12 I__7715 (
            .O(N__37508),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__7714 (
            .O(N__37503),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__7713 (
            .O(N__37498),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__7712 (
            .O(N__37495),
            .I(N__37492));
    LocalMux I__7711 (
            .O(N__37492),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__7710 (
            .O(N__37489),
            .I(N__37486));
    InMux I__7709 (
            .O(N__37486),
            .I(N__37483));
    LocalMux I__7708 (
            .O(N__37483),
            .I(N__37479));
    InMux I__7707 (
            .O(N__37482),
            .I(N__37476));
    Span4Mux_v I__7706 (
            .O(N__37479),
            .I(N__37472));
    LocalMux I__7705 (
            .O(N__37476),
            .I(N__37468));
    InMux I__7704 (
            .O(N__37475),
            .I(N__37465));
    Span4Mux_v I__7703 (
            .O(N__37472),
            .I(N__37462));
    InMux I__7702 (
            .O(N__37471),
            .I(N__37459));
    Span4Mux_v I__7701 (
            .O(N__37468),
            .I(N__37456));
    LocalMux I__7700 (
            .O(N__37465),
            .I(N__37453));
    Sp12to4 I__7699 (
            .O(N__37462),
            .I(N__37450));
    LocalMux I__7698 (
            .O(N__37459),
            .I(N__37447));
    Odrv4 I__7697 (
            .O(N__37456),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__7696 (
            .O(N__37453),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__7695 (
            .O(N__37450),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__7694 (
            .O(N__37447),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__7693 (
            .O(N__37438),
            .I(bfn_14_18_0_));
    InMux I__7692 (
            .O(N__37435),
            .I(N__37431));
    CascadeMux I__7691 (
            .O(N__37434),
            .I(N__37428));
    LocalMux I__7690 (
            .O(N__37431),
            .I(N__37424));
    InMux I__7689 (
            .O(N__37428),
            .I(N__37421));
    CascadeMux I__7688 (
            .O(N__37427),
            .I(N__37418));
    Span4Mux_v I__7687 (
            .O(N__37424),
            .I(N__37415));
    LocalMux I__7686 (
            .O(N__37421),
            .I(N__37411));
    InMux I__7685 (
            .O(N__37418),
            .I(N__37408));
    Span4Mux_h I__7684 (
            .O(N__37415),
            .I(N__37405));
    InMux I__7683 (
            .O(N__37414),
            .I(N__37402));
    Span4Mux_h I__7682 (
            .O(N__37411),
            .I(N__37397));
    LocalMux I__7681 (
            .O(N__37408),
            .I(N__37397));
    Span4Mux_h I__7680 (
            .O(N__37405),
            .I(N__37394));
    LocalMux I__7679 (
            .O(N__37402),
            .I(N__37391));
    Span4Mux_v I__7678 (
            .O(N__37397),
            .I(N__37388));
    Span4Mux_v I__7677 (
            .O(N__37394),
            .I(N__37383));
    Span4Mux_v I__7676 (
            .O(N__37391),
            .I(N__37383));
    Odrv4 I__7675 (
            .O(N__37388),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__7674 (
            .O(N__37383),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__7673 (
            .O(N__37378),
            .I(N__37375));
    InMux I__7672 (
            .O(N__37375),
            .I(N__37372));
    LocalMux I__7671 (
            .O(N__37372),
            .I(N__37369));
    Odrv12 I__7670 (
            .O(N__37369),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__7669 (
            .O(N__37366),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__7668 (
            .O(N__37363),
            .I(N__37360));
    LocalMux I__7667 (
            .O(N__37360),
            .I(N__37357));
    Span4Mux_h I__7666 (
            .O(N__37357),
            .I(N__37354));
    Odrv4 I__7665 (
            .O(N__37354),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__7664 (
            .O(N__37351),
            .I(N__37348));
    InMux I__7663 (
            .O(N__37348),
            .I(N__37345));
    LocalMux I__7662 (
            .O(N__37345),
            .I(N__37342));
    Span4Mux_v I__7661 (
            .O(N__37342),
            .I(N__37337));
    InMux I__7660 (
            .O(N__37341),
            .I(N__37334));
    InMux I__7659 (
            .O(N__37340),
            .I(N__37331));
    Span4Mux_h I__7658 (
            .O(N__37337),
            .I(N__37327));
    LocalMux I__7657 (
            .O(N__37334),
            .I(N__37324));
    LocalMux I__7656 (
            .O(N__37331),
            .I(N__37321));
    InMux I__7655 (
            .O(N__37330),
            .I(N__37318));
    Span4Mux_h I__7654 (
            .O(N__37327),
            .I(N__37313));
    Span4Mux_v I__7653 (
            .O(N__37324),
            .I(N__37313));
    Odrv4 I__7652 (
            .O(N__37321),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__7651 (
            .O(N__37318),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__7650 (
            .O(N__37313),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__7649 (
            .O(N__37306),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__7648 (
            .O(N__37303),
            .I(N__37300));
    LocalMux I__7647 (
            .O(N__37300),
            .I(N__37297));
    Odrv4 I__7646 (
            .O(N__37297),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__7645 (
            .O(N__37294),
            .I(N__37291));
    InMux I__7644 (
            .O(N__37291),
            .I(N__37288));
    LocalMux I__7643 (
            .O(N__37288),
            .I(N__37284));
    InMux I__7642 (
            .O(N__37287),
            .I(N__37280));
    Span4Mux_v I__7641 (
            .O(N__37284),
            .I(N__37277));
    InMux I__7640 (
            .O(N__37283),
            .I(N__37274));
    LocalMux I__7639 (
            .O(N__37280),
            .I(N__37271));
    Span4Mux_h I__7638 (
            .O(N__37277),
            .I(N__37268));
    LocalMux I__7637 (
            .O(N__37274),
            .I(N__37264));
    Span4Mux_h I__7636 (
            .O(N__37271),
            .I(N__37259));
    Span4Mux_h I__7635 (
            .O(N__37268),
            .I(N__37259));
    InMux I__7634 (
            .O(N__37267),
            .I(N__37256));
    Span4Mux_v I__7633 (
            .O(N__37264),
            .I(N__37253));
    Span4Mux_v I__7632 (
            .O(N__37259),
            .I(N__37248));
    LocalMux I__7631 (
            .O(N__37256),
            .I(N__37248));
    Odrv4 I__7630 (
            .O(N__37253),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__7629 (
            .O(N__37248),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__7628 (
            .O(N__37243),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__7627 (
            .O(N__37240),
            .I(N__37237));
    LocalMux I__7626 (
            .O(N__37237),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__7625 (
            .O(N__37234),
            .I(N__37231));
    InMux I__7624 (
            .O(N__37231),
            .I(N__37228));
    LocalMux I__7623 (
            .O(N__37228),
            .I(N__37225));
    Span4Mux_v I__7622 (
            .O(N__37225),
            .I(N__37220));
    InMux I__7621 (
            .O(N__37224),
            .I(N__37217));
    InMux I__7620 (
            .O(N__37223),
            .I(N__37214));
    Span4Mux_h I__7619 (
            .O(N__37220),
            .I(N__37211));
    LocalMux I__7618 (
            .O(N__37217),
            .I(N__37208));
    LocalMux I__7617 (
            .O(N__37214),
            .I(N__37204));
    Span4Mux_h I__7616 (
            .O(N__37211),
            .I(N__37201));
    Span4Mux_v I__7615 (
            .O(N__37208),
            .I(N__37198));
    InMux I__7614 (
            .O(N__37207),
            .I(N__37195));
    Span4Mux_v I__7613 (
            .O(N__37204),
            .I(N__37190));
    Span4Mux_h I__7612 (
            .O(N__37201),
            .I(N__37190));
    Odrv4 I__7611 (
            .O(N__37198),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__7610 (
            .O(N__37195),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__7609 (
            .O(N__37190),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__7608 (
            .O(N__37183),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__7607 (
            .O(N__37180),
            .I(N__37177));
    LocalMux I__7606 (
            .O(N__37177),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__7605 (
            .O(N__37174),
            .I(N__37171));
    InMux I__7604 (
            .O(N__37171),
            .I(N__37167));
    CascadeMux I__7603 (
            .O(N__37170),
            .I(N__37164));
    LocalMux I__7602 (
            .O(N__37167),
            .I(N__37160));
    InMux I__7601 (
            .O(N__37164),
            .I(N__37157));
    InMux I__7600 (
            .O(N__37163),
            .I(N__37154));
    Sp12to4 I__7599 (
            .O(N__37160),
            .I(N__37150));
    LocalMux I__7598 (
            .O(N__37157),
            .I(N__37145));
    LocalMux I__7597 (
            .O(N__37154),
            .I(N__37145));
    InMux I__7596 (
            .O(N__37153),
            .I(N__37142));
    Span12Mux_v I__7595 (
            .O(N__37150),
            .I(N__37139));
    Span4Mux_v I__7594 (
            .O(N__37145),
            .I(N__37136));
    LocalMux I__7593 (
            .O(N__37142),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv12 I__7592 (
            .O(N__37139),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__7591 (
            .O(N__37136),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__7590 (
            .O(N__37129),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__7589 (
            .O(N__37126),
            .I(N__37121));
    InMux I__7588 (
            .O(N__37125),
            .I(N__37116));
    InMux I__7587 (
            .O(N__37124),
            .I(N__37116));
    LocalMux I__7586 (
            .O(N__37121),
            .I(N__37110));
    LocalMux I__7585 (
            .O(N__37116),
            .I(N__37110));
    CascadeMux I__7584 (
            .O(N__37115),
            .I(N__37107));
    Sp12to4 I__7583 (
            .O(N__37110),
            .I(N__37104));
    InMux I__7582 (
            .O(N__37107),
            .I(N__37101));
    Span12Mux_v I__7581 (
            .O(N__37104),
            .I(N__37098));
    LocalMux I__7580 (
            .O(N__37101),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__7579 (
            .O(N__37098),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__7578 (
            .O(N__37093),
            .I(N__37090));
    LocalMux I__7577 (
            .O(N__37090),
            .I(N__37087));
    Odrv12 I__7576 (
            .O(N__37087),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__7575 (
            .O(N__37084),
            .I(N__37081));
    InMux I__7574 (
            .O(N__37081),
            .I(N__37077));
    InMux I__7573 (
            .O(N__37080),
            .I(N__37074));
    LocalMux I__7572 (
            .O(N__37077),
            .I(N__37071));
    LocalMux I__7571 (
            .O(N__37074),
            .I(N__37068));
    Sp12to4 I__7570 (
            .O(N__37071),
            .I(N__37065));
    Span4Mux_h I__7569 (
            .O(N__37068),
            .I(N__37061));
    Span12Mux_v I__7568 (
            .O(N__37065),
            .I(N__37058));
    InMux I__7567 (
            .O(N__37064),
            .I(N__37055));
    Sp12to4 I__7566 (
            .O(N__37061),
            .I(N__37050));
    Span12Mux_h I__7565 (
            .O(N__37058),
            .I(N__37050));
    LocalMux I__7564 (
            .O(N__37055),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv12 I__7563 (
            .O(N__37050),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__7562 (
            .O(N__37045),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__7561 (
            .O(N__37042),
            .I(N__37039));
    LocalMux I__7560 (
            .O(N__37039),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__7559 (
            .O(N__37036),
            .I(N__37032));
    InMux I__7558 (
            .O(N__37035),
            .I(N__37029));
    InMux I__7557 (
            .O(N__37032),
            .I(N__37026));
    LocalMux I__7556 (
            .O(N__37029),
            .I(N__37022));
    LocalMux I__7555 (
            .O(N__37026),
            .I(N__37019));
    InMux I__7554 (
            .O(N__37025),
            .I(N__37016));
    Span4Mux_v I__7553 (
            .O(N__37022),
            .I(N__37013));
    Span4Mux_v I__7552 (
            .O(N__37019),
            .I(N__37010));
    LocalMux I__7551 (
            .O(N__37016),
            .I(N__37007));
    Sp12to4 I__7550 (
            .O(N__37013),
            .I(N__37001));
    Sp12to4 I__7549 (
            .O(N__37010),
            .I(N__37001));
    Span4Mux_v I__7548 (
            .O(N__37007),
            .I(N__36998));
    InMux I__7547 (
            .O(N__37006),
            .I(N__36995));
    Span12Mux_h I__7546 (
            .O(N__37001),
            .I(N__36992));
    Odrv4 I__7545 (
            .O(N__36998),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__7544 (
            .O(N__36995),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__7543 (
            .O(N__36992),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__7542 (
            .O(N__36985),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__7541 (
            .O(N__36982),
            .I(N__36979));
    LocalMux I__7540 (
            .O(N__36979),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__7539 (
            .O(N__36976),
            .I(N__36972));
    InMux I__7538 (
            .O(N__36975),
            .I(N__36969));
    InMux I__7537 (
            .O(N__36972),
            .I(N__36966));
    LocalMux I__7536 (
            .O(N__36969),
            .I(N__36962));
    LocalMux I__7535 (
            .O(N__36966),
            .I(N__36959));
    InMux I__7534 (
            .O(N__36965),
            .I(N__36956));
    Span4Mux_v I__7533 (
            .O(N__36962),
            .I(N__36953));
    Span4Mux_v I__7532 (
            .O(N__36959),
            .I(N__36950));
    LocalMux I__7531 (
            .O(N__36956),
            .I(N__36947));
    Sp12to4 I__7530 (
            .O(N__36953),
            .I(N__36941));
    Sp12to4 I__7529 (
            .O(N__36950),
            .I(N__36941));
    Span4Mux_v I__7528 (
            .O(N__36947),
            .I(N__36938));
    InMux I__7527 (
            .O(N__36946),
            .I(N__36935));
    Span12Mux_h I__7526 (
            .O(N__36941),
            .I(N__36932));
    Odrv4 I__7525 (
            .O(N__36938),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__7524 (
            .O(N__36935),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__7523 (
            .O(N__36932),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__7522 (
            .O(N__36925),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__7521 (
            .O(N__36922),
            .I(N__36919));
    InMux I__7520 (
            .O(N__36919),
            .I(N__36916));
    LocalMux I__7519 (
            .O(N__36916),
            .I(N__36911));
    InMux I__7518 (
            .O(N__36915),
            .I(N__36907));
    InMux I__7517 (
            .O(N__36914),
            .I(N__36904));
    Span4Mux_v I__7516 (
            .O(N__36911),
            .I(N__36901));
    InMux I__7515 (
            .O(N__36910),
            .I(N__36898));
    LocalMux I__7514 (
            .O(N__36907),
            .I(N__36895));
    LocalMux I__7513 (
            .O(N__36904),
            .I(N__36892));
    Span4Mux_h I__7512 (
            .O(N__36901),
            .I(N__36889));
    LocalMux I__7511 (
            .O(N__36898),
            .I(N__36886));
    Span4Mux_h I__7510 (
            .O(N__36895),
            .I(N__36883));
    Span4Mux_h I__7509 (
            .O(N__36892),
            .I(N__36880));
    Sp12to4 I__7508 (
            .O(N__36889),
            .I(N__36877));
    Span4Mux_v I__7507 (
            .O(N__36886),
            .I(N__36874));
    Odrv4 I__7506 (
            .O(N__36883),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__7505 (
            .O(N__36880),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv12 I__7504 (
            .O(N__36877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__7503 (
            .O(N__36874),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__7502 (
            .O(N__36865),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__7501 (
            .O(N__36862),
            .I(N__36859));
    LocalMux I__7500 (
            .O(N__36859),
            .I(N__36856));
    Odrv4 I__7499 (
            .O(N__36856),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__7498 (
            .O(N__36853),
            .I(N__36850));
    InMux I__7497 (
            .O(N__36850),
            .I(N__36845));
    InMux I__7496 (
            .O(N__36849),
            .I(N__36842));
    CascadeMux I__7495 (
            .O(N__36848),
            .I(N__36839));
    LocalMux I__7494 (
            .O(N__36845),
            .I(N__36836));
    LocalMux I__7493 (
            .O(N__36842),
            .I(N__36833));
    InMux I__7492 (
            .O(N__36839),
            .I(N__36830));
    Span4Mux_v I__7491 (
            .O(N__36836),
            .I(N__36827));
    Span4Mux_h I__7490 (
            .O(N__36833),
            .I(N__36824));
    LocalMux I__7489 (
            .O(N__36830),
            .I(N__36821));
    Span4Mux_v I__7488 (
            .O(N__36827),
            .I(N__36817));
    Span4Mux_v I__7487 (
            .O(N__36824),
            .I(N__36814));
    Span4Mux_v I__7486 (
            .O(N__36821),
            .I(N__36811));
    InMux I__7485 (
            .O(N__36820),
            .I(N__36808));
    Sp12to4 I__7484 (
            .O(N__36817),
            .I(N__36805));
    Odrv4 I__7483 (
            .O(N__36814),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__7482 (
            .O(N__36811),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__7481 (
            .O(N__36808),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv12 I__7480 (
            .O(N__36805),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__7479 (
            .O(N__36796),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__7478 (
            .O(N__36793),
            .I(N__36787));
    InMux I__7477 (
            .O(N__36792),
            .I(N__36787));
    LocalMux I__7476 (
            .O(N__36787),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    CascadeMux I__7475 (
            .O(N__36784),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ));
    InMux I__7474 (
            .O(N__36781),
            .I(N__36775));
    InMux I__7473 (
            .O(N__36780),
            .I(N__36775));
    LocalMux I__7472 (
            .O(N__36775),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__7471 (
            .O(N__36772),
            .I(N__36768));
    InMux I__7470 (
            .O(N__36771),
            .I(N__36764));
    LocalMux I__7469 (
            .O(N__36768),
            .I(N__36761));
    InMux I__7468 (
            .O(N__36767),
            .I(N__36758));
    LocalMux I__7467 (
            .O(N__36764),
            .I(N__36755));
    Span4Mux_v I__7466 (
            .O(N__36761),
            .I(N__36750));
    LocalMux I__7465 (
            .O(N__36758),
            .I(N__36750));
    Span4Mux_h I__7464 (
            .O(N__36755),
            .I(N__36747));
    Odrv4 I__7463 (
            .O(N__36750),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7462 (
            .O(N__36747),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__7461 (
            .O(N__36742),
            .I(N__36738));
    InMux I__7460 (
            .O(N__36741),
            .I(N__36735));
    LocalMux I__7459 (
            .O(N__36738),
            .I(N__36732));
    LocalMux I__7458 (
            .O(N__36735),
            .I(N__36729));
    Span4Mux_s3_h I__7457 (
            .O(N__36732),
            .I(N__36726));
    Span4Mux_h I__7456 (
            .O(N__36729),
            .I(N__36723));
    Span4Mux_h I__7455 (
            .O(N__36726),
            .I(N__36720));
    Odrv4 I__7454 (
            .O(N__36723),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__7453 (
            .O(N__36720),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__7452 (
            .O(N__36715),
            .I(N__36711));
    InMux I__7451 (
            .O(N__36714),
            .I(N__36708));
    LocalMux I__7450 (
            .O(N__36711),
            .I(N__36705));
    LocalMux I__7449 (
            .O(N__36708),
            .I(N__36702));
    Span4Mux_h I__7448 (
            .O(N__36705),
            .I(N__36699));
    Span4Mux_s3_h I__7447 (
            .O(N__36702),
            .I(N__36696));
    Span4Mux_h I__7446 (
            .O(N__36699),
            .I(N__36693));
    Span4Mux_h I__7445 (
            .O(N__36696),
            .I(N__36690));
    Odrv4 I__7444 (
            .O(N__36693),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__7443 (
            .O(N__36690),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__7442 (
            .O(N__36685),
            .I(N__36681));
    InMux I__7441 (
            .O(N__36684),
            .I(N__36678));
    LocalMux I__7440 (
            .O(N__36681),
            .I(N__36675));
    LocalMux I__7439 (
            .O(N__36678),
            .I(N__36672));
    Span4Mux_v I__7438 (
            .O(N__36675),
            .I(N__36669));
    Span4Mux_v I__7437 (
            .O(N__36672),
            .I(N__36666));
    Sp12to4 I__7436 (
            .O(N__36669),
            .I(N__36663));
    Span4Mux_h I__7435 (
            .O(N__36666),
            .I(N__36660));
    Odrv12 I__7434 (
            .O(N__36663),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__7433 (
            .O(N__36660),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__7432 (
            .O(N__36655),
            .I(N__36649));
    InMux I__7431 (
            .O(N__36654),
            .I(N__36649));
    LocalMux I__7430 (
            .O(N__36649),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    InMux I__7429 (
            .O(N__36646),
            .I(N__36642));
    InMux I__7428 (
            .O(N__36645),
            .I(N__36639));
    LocalMux I__7427 (
            .O(N__36642),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    LocalMux I__7426 (
            .O(N__36639),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__7425 (
            .O(N__36634),
            .I(N__36630));
    InMux I__7424 (
            .O(N__36633),
            .I(N__36627));
    LocalMux I__7423 (
            .O(N__36630),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    LocalMux I__7422 (
            .O(N__36627),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    CascadeMux I__7421 (
            .O(N__36622),
            .I(N__36619));
    InMux I__7420 (
            .O(N__36619),
            .I(N__36616));
    LocalMux I__7419 (
            .O(N__36616),
            .I(N__36613));
    Odrv4 I__7418 (
            .O(N__36613),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__7417 (
            .O(N__36610),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__7416 (
            .O(N__36607),
            .I(N__36604));
    LocalMux I__7415 (
            .O(N__36604),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ));
    CascadeMux I__7414 (
            .O(N__36601),
            .I(N__36597));
    CascadeMux I__7413 (
            .O(N__36600),
            .I(N__36594));
    InMux I__7412 (
            .O(N__36597),
            .I(N__36589));
    InMux I__7411 (
            .O(N__36594),
            .I(N__36589));
    LocalMux I__7410 (
            .O(N__36589),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    CascadeMux I__7409 (
            .O(N__36586),
            .I(N__36583));
    InMux I__7408 (
            .O(N__36583),
            .I(N__36578));
    InMux I__7407 (
            .O(N__36582),
            .I(N__36575));
    InMux I__7406 (
            .O(N__36581),
            .I(N__36572));
    LocalMux I__7405 (
            .O(N__36578),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__7404 (
            .O(N__36575),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__7403 (
            .O(N__36572),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__7402 (
            .O(N__36565),
            .I(bfn_14_10_0_));
    CascadeMux I__7401 (
            .O(N__36562),
            .I(N__36559));
    InMux I__7400 (
            .O(N__36559),
            .I(N__36554));
    InMux I__7399 (
            .O(N__36558),
            .I(N__36551));
    InMux I__7398 (
            .O(N__36557),
            .I(N__36548));
    LocalMux I__7397 (
            .O(N__36554),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__7396 (
            .O(N__36551),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__7395 (
            .O(N__36548),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__7394 (
            .O(N__36541),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7393 (
            .O(N__36538),
            .I(N__36534));
    InMux I__7392 (
            .O(N__36537),
            .I(N__36531));
    LocalMux I__7391 (
            .O(N__36534),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__7390 (
            .O(N__36531),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__7389 (
            .O(N__36526),
            .I(N__36523));
    InMux I__7388 (
            .O(N__36523),
            .I(N__36518));
    InMux I__7387 (
            .O(N__36522),
            .I(N__36515));
    InMux I__7386 (
            .O(N__36521),
            .I(N__36512));
    LocalMux I__7385 (
            .O(N__36518),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__7384 (
            .O(N__36515),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__7383 (
            .O(N__36512),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__7382 (
            .O(N__36505),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__7381 (
            .O(N__36502),
            .I(N__36498));
    InMux I__7380 (
            .O(N__36501),
            .I(N__36495));
    LocalMux I__7379 (
            .O(N__36498),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__7378 (
            .O(N__36495),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__7377 (
            .O(N__36490),
            .I(N__36487));
    InMux I__7376 (
            .O(N__36487),
            .I(N__36482));
    InMux I__7375 (
            .O(N__36486),
            .I(N__36479));
    InMux I__7374 (
            .O(N__36485),
            .I(N__36476));
    LocalMux I__7373 (
            .O(N__36482),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__7372 (
            .O(N__36479),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__7371 (
            .O(N__36476),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__7370 (
            .O(N__36469),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7369 (
            .O(N__36466),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__7368 (
            .O(N__36463),
            .I(N__36457));
    CEMux I__7367 (
            .O(N__36462),
            .I(N__36454));
    CEMux I__7366 (
            .O(N__36461),
            .I(N__36451));
    CEMux I__7365 (
            .O(N__36460),
            .I(N__36448));
    LocalMux I__7364 (
            .O(N__36457),
            .I(N__36444));
    LocalMux I__7363 (
            .O(N__36454),
            .I(N__36441));
    LocalMux I__7362 (
            .O(N__36451),
            .I(N__36438));
    LocalMux I__7361 (
            .O(N__36448),
            .I(N__36435));
    CEMux I__7360 (
            .O(N__36447),
            .I(N__36432));
    Span4Mux_h I__7359 (
            .O(N__36444),
            .I(N__36429));
    Span4Mux_h I__7358 (
            .O(N__36441),
            .I(N__36426));
    Span4Mux_h I__7357 (
            .O(N__36438),
            .I(N__36423));
    Span4Mux_h I__7356 (
            .O(N__36435),
            .I(N__36420));
    LocalMux I__7355 (
            .O(N__36432),
            .I(N__36417));
    Odrv4 I__7354 (
            .O(N__36429),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__7353 (
            .O(N__36426),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__7352 (
            .O(N__36423),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__7351 (
            .O(N__36420),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv12 I__7350 (
            .O(N__36417),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    CascadeMux I__7349 (
            .O(N__36406),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_));
    CascadeMux I__7348 (
            .O(N__36403),
            .I(N__36400));
    InMux I__7347 (
            .O(N__36400),
            .I(N__36394));
    InMux I__7346 (
            .O(N__36399),
            .I(N__36394));
    LocalMux I__7345 (
            .O(N__36394),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    CascadeMux I__7344 (
            .O(N__36391),
            .I(N__36388));
    InMux I__7343 (
            .O(N__36388),
            .I(N__36383));
    InMux I__7342 (
            .O(N__36387),
            .I(N__36380));
    InMux I__7341 (
            .O(N__36386),
            .I(N__36377));
    LocalMux I__7340 (
            .O(N__36383),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__7339 (
            .O(N__36380),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__7338 (
            .O(N__36377),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__7337 (
            .O(N__36370),
            .I(bfn_14_9_0_));
    CascadeMux I__7336 (
            .O(N__36367),
            .I(N__36364));
    InMux I__7335 (
            .O(N__36364),
            .I(N__36359));
    InMux I__7334 (
            .O(N__36363),
            .I(N__36356));
    InMux I__7333 (
            .O(N__36362),
            .I(N__36353));
    LocalMux I__7332 (
            .O(N__36359),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__7331 (
            .O(N__36356),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__7330 (
            .O(N__36353),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__7329 (
            .O(N__36346),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__7328 (
            .O(N__36343),
            .I(N__36338));
    InMux I__7327 (
            .O(N__36342),
            .I(N__36333));
    InMux I__7326 (
            .O(N__36341),
            .I(N__36333));
    LocalMux I__7325 (
            .O(N__36338),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__7324 (
            .O(N__36333),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__7323 (
            .O(N__36328),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__7322 (
            .O(N__36325),
            .I(N__36322));
    InMux I__7321 (
            .O(N__36322),
            .I(N__36317));
    InMux I__7320 (
            .O(N__36321),
            .I(N__36314));
    InMux I__7319 (
            .O(N__36320),
            .I(N__36311));
    LocalMux I__7318 (
            .O(N__36317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__7317 (
            .O(N__36314),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__7316 (
            .O(N__36311),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__7315 (
            .O(N__36304),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__7314 (
            .O(N__36301),
            .I(N__36296));
    CascadeMux I__7313 (
            .O(N__36300),
            .I(N__36293));
    InMux I__7312 (
            .O(N__36299),
            .I(N__36290));
    InMux I__7311 (
            .O(N__36296),
            .I(N__36285));
    InMux I__7310 (
            .O(N__36293),
            .I(N__36285));
    LocalMux I__7309 (
            .O(N__36290),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__7308 (
            .O(N__36285),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__7307 (
            .O(N__36280),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__7306 (
            .O(N__36277),
            .I(N__36274));
    InMux I__7305 (
            .O(N__36274),
            .I(N__36269));
    InMux I__7304 (
            .O(N__36273),
            .I(N__36266));
    InMux I__7303 (
            .O(N__36272),
            .I(N__36263));
    LocalMux I__7302 (
            .O(N__36269),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__7301 (
            .O(N__36266),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__7300 (
            .O(N__36263),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__7299 (
            .O(N__36256),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__7298 (
            .O(N__36253),
            .I(N__36250));
    InMux I__7297 (
            .O(N__36250),
            .I(N__36245));
    InMux I__7296 (
            .O(N__36249),
            .I(N__36242));
    InMux I__7295 (
            .O(N__36248),
            .I(N__36239));
    LocalMux I__7294 (
            .O(N__36245),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__7293 (
            .O(N__36242),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__7292 (
            .O(N__36239),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__7291 (
            .O(N__36232),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7290 (
            .O(N__36229),
            .I(N__36226));
    InMux I__7289 (
            .O(N__36226),
            .I(N__36221));
    InMux I__7288 (
            .O(N__36225),
            .I(N__36218));
    InMux I__7287 (
            .O(N__36224),
            .I(N__36215));
    LocalMux I__7286 (
            .O(N__36221),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__7285 (
            .O(N__36218),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__7284 (
            .O(N__36215),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__7283 (
            .O(N__36208),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__7282 (
            .O(N__36205),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7281 (
            .O(N__36202),
            .I(N__36199));
    InMux I__7280 (
            .O(N__36199),
            .I(N__36194));
    InMux I__7279 (
            .O(N__36198),
            .I(N__36191));
    InMux I__7278 (
            .O(N__36197),
            .I(N__36188));
    LocalMux I__7277 (
            .O(N__36194),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__7276 (
            .O(N__36191),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__7275 (
            .O(N__36188),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__7274 (
            .O(N__36181),
            .I(bfn_14_8_0_));
    CascadeMux I__7273 (
            .O(N__36178),
            .I(N__36175));
    InMux I__7272 (
            .O(N__36175),
            .I(N__36170));
    InMux I__7271 (
            .O(N__36174),
            .I(N__36167));
    InMux I__7270 (
            .O(N__36173),
            .I(N__36164));
    LocalMux I__7269 (
            .O(N__36170),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__7268 (
            .O(N__36167),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__7267 (
            .O(N__36164),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__7266 (
            .O(N__36157),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7265 (
            .O(N__36154),
            .I(N__36151));
    InMux I__7264 (
            .O(N__36151),
            .I(N__36146));
    InMux I__7263 (
            .O(N__36150),
            .I(N__36143));
    InMux I__7262 (
            .O(N__36149),
            .I(N__36140));
    LocalMux I__7261 (
            .O(N__36146),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__7260 (
            .O(N__36143),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__7259 (
            .O(N__36140),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__7258 (
            .O(N__36133),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__7257 (
            .O(N__36130),
            .I(N__36127));
    InMux I__7256 (
            .O(N__36127),
            .I(N__36122));
    InMux I__7255 (
            .O(N__36126),
            .I(N__36119));
    InMux I__7254 (
            .O(N__36125),
            .I(N__36116));
    LocalMux I__7253 (
            .O(N__36122),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__7252 (
            .O(N__36119),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__7251 (
            .O(N__36116),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__7250 (
            .O(N__36109),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__7249 (
            .O(N__36106),
            .I(N__36103));
    InMux I__7248 (
            .O(N__36103),
            .I(N__36098));
    InMux I__7247 (
            .O(N__36102),
            .I(N__36095));
    InMux I__7246 (
            .O(N__36101),
            .I(N__36092));
    LocalMux I__7245 (
            .O(N__36098),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__7244 (
            .O(N__36095),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__7243 (
            .O(N__36092),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__7242 (
            .O(N__36085),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__7241 (
            .O(N__36082),
            .I(N__36079));
    InMux I__7240 (
            .O(N__36079),
            .I(N__36074));
    InMux I__7239 (
            .O(N__36078),
            .I(N__36071));
    InMux I__7238 (
            .O(N__36077),
            .I(N__36068));
    LocalMux I__7237 (
            .O(N__36074),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__7236 (
            .O(N__36071),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__7235 (
            .O(N__36068),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__7234 (
            .O(N__36061),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7233 (
            .O(N__36058),
            .I(N__36055));
    InMux I__7232 (
            .O(N__36055),
            .I(N__36050));
    InMux I__7231 (
            .O(N__36054),
            .I(N__36047));
    InMux I__7230 (
            .O(N__36053),
            .I(N__36044));
    LocalMux I__7229 (
            .O(N__36050),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__7228 (
            .O(N__36047),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__7227 (
            .O(N__36044),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__7226 (
            .O(N__36037),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__7225 (
            .O(N__36034),
            .I(N__36031));
    InMux I__7224 (
            .O(N__36031),
            .I(N__36026));
    InMux I__7223 (
            .O(N__36030),
            .I(N__36023));
    InMux I__7222 (
            .O(N__36029),
            .I(N__36020));
    LocalMux I__7221 (
            .O(N__36026),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__7220 (
            .O(N__36023),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__7219 (
            .O(N__36020),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__7218 (
            .O(N__36013),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__7217 (
            .O(N__36010),
            .I(N__36006));
    InMux I__7216 (
            .O(N__36009),
            .I(N__36002));
    InMux I__7215 (
            .O(N__36006),
            .I(N__35999));
    InMux I__7214 (
            .O(N__36005),
            .I(N__35996));
    LocalMux I__7213 (
            .O(N__36002),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__7212 (
            .O(N__35999),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__7211 (
            .O(N__35996),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__7210 (
            .O(N__35989),
            .I(N__35985));
    InMux I__7209 (
            .O(N__35988),
            .I(N__35981));
    InMux I__7208 (
            .O(N__35985),
            .I(N__35978));
    InMux I__7207 (
            .O(N__35984),
            .I(N__35975));
    LocalMux I__7206 (
            .O(N__35981),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__7205 (
            .O(N__35978),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__7204 (
            .O(N__35975),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__7203 (
            .O(N__35968),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__7202 (
            .O(N__35965),
            .I(N__35962));
    InMux I__7201 (
            .O(N__35962),
            .I(N__35957));
    InMux I__7200 (
            .O(N__35961),
            .I(N__35954));
    InMux I__7199 (
            .O(N__35960),
            .I(N__35951));
    LocalMux I__7198 (
            .O(N__35957),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__7197 (
            .O(N__35954),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__7196 (
            .O(N__35951),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__7195 (
            .O(N__35944),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__7194 (
            .O(N__35941),
            .I(N__35938));
    InMux I__7193 (
            .O(N__35938),
            .I(N__35933));
    InMux I__7192 (
            .O(N__35937),
            .I(N__35930));
    InMux I__7191 (
            .O(N__35936),
            .I(N__35927));
    LocalMux I__7190 (
            .O(N__35933),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__7189 (
            .O(N__35930),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__7188 (
            .O(N__35927),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__7187 (
            .O(N__35920),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__7186 (
            .O(N__35917),
            .I(N__35914));
    InMux I__7185 (
            .O(N__35914),
            .I(N__35909));
    InMux I__7184 (
            .O(N__35913),
            .I(N__35906));
    InMux I__7183 (
            .O(N__35912),
            .I(N__35903));
    LocalMux I__7182 (
            .O(N__35909),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__7181 (
            .O(N__35906),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__7180 (
            .O(N__35903),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__7179 (
            .O(N__35896),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__7178 (
            .O(N__35893),
            .I(N__35890));
    InMux I__7177 (
            .O(N__35890),
            .I(N__35885));
    InMux I__7176 (
            .O(N__35889),
            .I(N__35882));
    InMux I__7175 (
            .O(N__35888),
            .I(N__35879));
    LocalMux I__7174 (
            .O(N__35885),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__7173 (
            .O(N__35882),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__7172 (
            .O(N__35879),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__7171 (
            .O(N__35872),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7170 (
            .O(N__35869),
            .I(N__35866));
    InMux I__7169 (
            .O(N__35866),
            .I(N__35861));
    InMux I__7168 (
            .O(N__35865),
            .I(N__35858));
    InMux I__7167 (
            .O(N__35864),
            .I(N__35855));
    LocalMux I__7166 (
            .O(N__35861),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__7165 (
            .O(N__35858),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__7164 (
            .O(N__35855),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__7163 (
            .O(N__35848),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7162 (
            .O(N__35845),
            .I(N__35842));
    InMux I__7161 (
            .O(N__35842),
            .I(N__35837));
    InMux I__7160 (
            .O(N__35841),
            .I(N__35834));
    InMux I__7159 (
            .O(N__35840),
            .I(N__35831));
    LocalMux I__7158 (
            .O(N__35837),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__7157 (
            .O(N__35834),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__7156 (
            .O(N__35831),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__7155 (
            .O(N__35824),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__7154 (
            .O(N__35821),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__7153 (
            .O(N__35818),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__7152 (
            .O(N__35815),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__7151 (
            .O(N__35812),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__7150 (
            .O(N__35809),
            .I(bfn_13_27_0_));
    InMux I__7149 (
            .O(N__35806),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    CascadeMux I__7148 (
            .O(N__35803),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ));
    CascadeMux I__7147 (
            .O(N__35800),
            .I(N__35797));
    InMux I__7146 (
            .O(N__35797),
            .I(N__35794));
    LocalMux I__7145 (
            .O(N__35794),
            .I(N__35791));
    Odrv4 I__7144 (
            .O(N__35791),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__7143 (
            .O(N__35788),
            .I(N__35783));
    InMux I__7142 (
            .O(N__35787),
            .I(N__35780));
    InMux I__7141 (
            .O(N__35786),
            .I(N__35777));
    LocalMux I__7140 (
            .O(N__35783),
            .I(N__35774));
    LocalMux I__7139 (
            .O(N__35780),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__7138 (
            .O(N__35777),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__7137 (
            .O(N__35774),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__7136 (
            .O(N__35767),
            .I(N__35764));
    LocalMux I__7135 (
            .O(N__35764),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__7134 (
            .O(N__35761),
            .I(N__35756));
    InMux I__7133 (
            .O(N__35760),
            .I(N__35753));
    InMux I__7132 (
            .O(N__35759),
            .I(N__35750));
    LocalMux I__7131 (
            .O(N__35756),
            .I(N__35747));
    LocalMux I__7130 (
            .O(N__35753),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__7129 (
            .O(N__35750),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__7128 (
            .O(N__35747),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__7127 (
            .O(N__35740),
            .I(N__35737));
    LocalMux I__7126 (
            .O(N__35737),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__7125 (
            .O(N__35734),
            .I(N__35729));
    InMux I__7124 (
            .O(N__35733),
            .I(N__35726));
    InMux I__7123 (
            .O(N__35732),
            .I(N__35723));
    LocalMux I__7122 (
            .O(N__35729),
            .I(N__35718));
    LocalMux I__7121 (
            .O(N__35726),
            .I(N__35718));
    LocalMux I__7120 (
            .O(N__35723),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__7119 (
            .O(N__35718),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__7118 (
            .O(N__35713),
            .I(N__35710));
    LocalMux I__7117 (
            .O(N__35710),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__7116 (
            .O(N__35707),
            .I(N__35702));
    InMux I__7115 (
            .O(N__35706),
            .I(N__35699));
    InMux I__7114 (
            .O(N__35705),
            .I(N__35696));
    LocalMux I__7113 (
            .O(N__35702),
            .I(N__35693));
    LocalMux I__7112 (
            .O(N__35699),
            .I(N__35690));
    LocalMux I__7111 (
            .O(N__35696),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__7110 (
            .O(N__35693),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__7109 (
            .O(N__35690),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__7108 (
            .O(N__35683),
            .I(N__35680));
    LocalMux I__7107 (
            .O(N__35680),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__7106 (
            .O(N__35677),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__7105 (
            .O(N__35674),
            .I(N__35671));
    LocalMux I__7104 (
            .O(N__35671),
            .I(N__35668));
    IoSpan4Mux I__7103 (
            .O(N__35668),
            .I(N__35665));
    Sp12to4 I__7102 (
            .O(N__35665),
            .I(N__35662));
    Span12Mux_s10_v I__7101 (
            .O(N__35662),
            .I(N__35659));
    Span12Mux_v I__7100 (
            .O(N__35659),
            .I(N__35656));
    Span12Mux_h I__7099 (
            .O(N__35656),
            .I(N__35653));
    Odrv12 I__7098 (
            .O(N__35653),
            .I(pwm_output_c));
    InMux I__7097 (
            .O(N__35650),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__7096 (
            .O(N__35647),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__7095 (
            .O(N__35644),
            .I(N__35640));
    InMux I__7094 (
            .O(N__35643),
            .I(N__35637));
    LocalMux I__7093 (
            .O(N__35640),
            .I(N__35634));
    LocalMux I__7092 (
            .O(N__35637),
            .I(N__35631));
    Span4Mux_s3_h I__7091 (
            .O(N__35634),
            .I(N__35628));
    Span4Mux_h I__7090 (
            .O(N__35631),
            .I(N__35625));
    Span4Mux_h I__7089 (
            .O(N__35628),
            .I(N__35622));
    Span4Mux_h I__7088 (
            .O(N__35625),
            .I(N__35619));
    Sp12to4 I__7087 (
            .O(N__35622),
            .I(N__35616));
    Odrv4 I__7086 (
            .O(N__35619),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv12 I__7085 (
            .O(N__35616),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__7084 (
            .O(N__35611),
            .I(N__35596));
    InMux I__7083 (
            .O(N__35610),
            .I(N__35596));
    InMux I__7082 (
            .O(N__35609),
            .I(N__35584));
    InMux I__7081 (
            .O(N__35608),
            .I(N__35584));
    InMux I__7080 (
            .O(N__35607),
            .I(N__35584));
    InMux I__7079 (
            .O(N__35606),
            .I(N__35584));
    InMux I__7078 (
            .O(N__35605),
            .I(N__35584));
    InMux I__7077 (
            .O(N__35604),
            .I(N__35557));
    InMux I__7076 (
            .O(N__35603),
            .I(N__35557));
    InMux I__7075 (
            .O(N__35602),
            .I(N__35554));
    InMux I__7074 (
            .O(N__35601),
            .I(N__35548));
    LocalMux I__7073 (
            .O(N__35596),
            .I(N__35545));
    InMux I__7072 (
            .O(N__35595),
            .I(N__35531));
    LocalMux I__7071 (
            .O(N__35584),
            .I(N__35528));
    InMux I__7070 (
            .O(N__35583),
            .I(N__35525));
    InMux I__7069 (
            .O(N__35582),
            .I(N__35520));
    InMux I__7068 (
            .O(N__35581),
            .I(N__35520));
    InMux I__7067 (
            .O(N__35580),
            .I(N__35513));
    InMux I__7066 (
            .O(N__35579),
            .I(N__35513));
    InMux I__7065 (
            .O(N__35578),
            .I(N__35513));
    InMux I__7064 (
            .O(N__35577),
            .I(N__35502));
    InMux I__7063 (
            .O(N__35576),
            .I(N__35502));
    InMux I__7062 (
            .O(N__35575),
            .I(N__35502));
    InMux I__7061 (
            .O(N__35574),
            .I(N__35502));
    InMux I__7060 (
            .O(N__35573),
            .I(N__35502));
    InMux I__7059 (
            .O(N__35572),
            .I(N__35493));
    InMux I__7058 (
            .O(N__35571),
            .I(N__35486));
    InMux I__7057 (
            .O(N__35570),
            .I(N__35486));
    InMux I__7056 (
            .O(N__35569),
            .I(N__35486));
    InMux I__7055 (
            .O(N__35568),
            .I(N__35471));
    InMux I__7054 (
            .O(N__35567),
            .I(N__35471));
    InMux I__7053 (
            .O(N__35566),
            .I(N__35471));
    InMux I__7052 (
            .O(N__35565),
            .I(N__35471));
    InMux I__7051 (
            .O(N__35564),
            .I(N__35471));
    InMux I__7050 (
            .O(N__35563),
            .I(N__35471));
    InMux I__7049 (
            .O(N__35562),
            .I(N__35471));
    LocalMux I__7048 (
            .O(N__35557),
            .I(N__35468));
    LocalMux I__7047 (
            .O(N__35554),
            .I(N__35465));
    InMux I__7046 (
            .O(N__35553),
            .I(N__35460));
    InMux I__7045 (
            .O(N__35552),
            .I(N__35460));
    InMux I__7044 (
            .O(N__35551),
            .I(N__35457));
    LocalMux I__7043 (
            .O(N__35548),
            .I(N__35444));
    Span4Mux_v I__7042 (
            .O(N__35545),
            .I(N__35444));
    InMux I__7041 (
            .O(N__35544),
            .I(N__35431));
    InMux I__7040 (
            .O(N__35543),
            .I(N__35431));
    InMux I__7039 (
            .O(N__35542),
            .I(N__35431));
    InMux I__7038 (
            .O(N__35541),
            .I(N__35431));
    InMux I__7037 (
            .O(N__35540),
            .I(N__35431));
    InMux I__7036 (
            .O(N__35539),
            .I(N__35431));
    InMux I__7035 (
            .O(N__35538),
            .I(N__35415));
    InMux I__7034 (
            .O(N__35537),
            .I(N__35415));
    InMux I__7033 (
            .O(N__35536),
            .I(N__35415));
    InMux I__7032 (
            .O(N__35535),
            .I(N__35412));
    InMux I__7031 (
            .O(N__35534),
            .I(N__35409));
    LocalMux I__7030 (
            .O(N__35531),
            .I(N__35396));
    Span4Mux_v I__7029 (
            .O(N__35528),
            .I(N__35396));
    LocalMux I__7028 (
            .O(N__35525),
            .I(N__35396));
    LocalMux I__7027 (
            .O(N__35520),
            .I(N__35396));
    LocalMux I__7026 (
            .O(N__35513),
            .I(N__35396));
    LocalMux I__7025 (
            .O(N__35502),
            .I(N__35396));
    InMux I__7024 (
            .O(N__35501),
            .I(N__35383));
    InMux I__7023 (
            .O(N__35500),
            .I(N__35383));
    InMux I__7022 (
            .O(N__35499),
            .I(N__35383));
    InMux I__7021 (
            .O(N__35498),
            .I(N__35383));
    InMux I__7020 (
            .O(N__35497),
            .I(N__35383));
    InMux I__7019 (
            .O(N__35496),
            .I(N__35383));
    LocalMux I__7018 (
            .O(N__35493),
            .I(N__35374));
    LocalMux I__7017 (
            .O(N__35486),
            .I(N__35374));
    LocalMux I__7016 (
            .O(N__35471),
            .I(N__35374));
    Span4Mux_h I__7015 (
            .O(N__35468),
            .I(N__35374));
    Span4Mux_h I__7014 (
            .O(N__35465),
            .I(N__35369));
    LocalMux I__7013 (
            .O(N__35460),
            .I(N__35369));
    LocalMux I__7012 (
            .O(N__35457),
            .I(N__35366));
    InMux I__7011 (
            .O(N__35456),
            .I(N__35349));
    InMux I__7010 (
            .O(N__35455),
            .I(N__35349));
    InMux I__7009 (
            .O(N__35454),
            .I(N__35349));
    InMux I__7008 (
            .O(N__35453),
            .I(N__35349));
    InMux I__7007 (
            .O(N__35452),
            .I(N__35349));
    InMux I__7006 (
            .O(N__35451),
            .I(N__35349));
    InMux I__7005 (
            .O(N__35450),
            .I(N__35349));
    InMux I__7004 (
            .O(N__35449),
            .I(N__35349));
    Span4Mux_v I__7003 (
            .O(N__35444),
            .I(N__35344));
    LocalMux I__7002 (
            .O(N__35431),
            .I(N__35344));
    InMux I__7001 (
            .O(N__35430),
            .I(N__35331));
    InMux I__7000 (
            .O(N__35429),
            .I(N__35331));
    InMux I__6999 (
            .O(N__35428),
            .I(N__35331));
    InMux I__6998 (
            .O(N__35427),
            .I(N__35331));
    InMux I__6997 (
            .O(N__35426),
            .I(N__35331));
    InMux I__6996 (
            .O(N__35425),
            .I(N__35331));
    InMux I__6995 (
            .O(N__35424),
            .I(N__35324));
    InMux I__6994 (
            .O(N__35423),
            .I(N__35324));
    InMux I__6993 (
            .O(N__35422),
            .I(N__35324));
    LocalMux I__6992 (
            .O(N__35415),
            .I(N__35321));
    LocalMux I__6991 (
            .O(N__35412),
            .I(N__35314));
    LocalMux I__6990 (
            .O(N__35409),
            .I(N__35314));
    Span4Mux_v I__6989 (
            .O(N__35396),
            .I(N__35314));
    LocalMux I__6988 (
            .O(N__35383),
            .I(N__35307));
    Span4Mux_v I__6987 (
            .O(N__35374),
            .I(N__35307));
    Span4Mux_h I__6986 (
            .O(N__35369),
            .I(N__35307));
    Odrv12 I__6985 (
            .O(N__35366),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6984 (
            .O(N__35349),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6983 (
            .O(N__35344),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6982 (
            .O(N__35331),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6981 (
            .O(N__35324),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__6980 (
            .O(N__35321),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6979 (
            .O(N__35314),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6978 (
            .O(N__35307),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__6977 (
            .O(N__35290),
            .I(N__35287));
    InMux I__6976 (
            .O(N__35287),
            .I(N__35284));
    LocalMux I__6975 (
            .O(N__35284),
            .I(N__35280));
    InMux I__6974 (
            .O(N__35283),
            .I(N__35276));
    Span4Mux_h I__6973 (
            .O(N__35280),
            .I(N__35273));
    InMux I__6972 (
            .O(N__35279),
            .I(N__35270));
    LocalMux I__6971 (
            .O(N__35276),
            .I(N__35267));
    Span4Mux_v I__6970 (
            .O(N__35273),
            .I(N__35263));
    LocalMux I__6969 (
            .O(N__35270),
            .I(N__35260));
    Span4Mux_h I__6968 (
            .O(N__35267),
            .I(N__35257));
    InMux I__6967 (
            .O(N__35266),
            .I(N__35254));
    Odrv4 I__6966 (
            .O(N__35263),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv12 I__6965 (
            .O(N__35260),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__6964 (
            .O(N__35257),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__6963 (
            .O(N__35254),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__6962 (
            .O(N__35245),
            .I(N__35210));
    InMux I__6961 (
            .O(N__35244),
            .I(N__35210));
    InMux I__6960 (
            .O(N__35243),
            .I(N__35199));
    InMux I__6959 (
            .O(N__35242),
            .I(N__35199));
    InMux I__6958 (
            .O(N__35241),
            .I(N__35199));
    InMux I__6957 (
            .O(N__35240),
            .I(N__35199));
    InMux I__6956 (
            .O(N__35239),
            .I(N__35199));
    CascadeMux I__6955 (
            .O(N__35238),
            .I(N__35194));
    CascadeMux I__6954 (
            .O(N__35237),
            .I(N__35189));
    InMux I__6953 (
            .O(N__35236),
            .I(N__35181));
    CascadeMux I__6952 (
            .O(N__35235),
            .I(N__35178));
    CascadeMux I__6951 (
            .O(N__35234),
            .I(N__35172));
    CascadeMux I__6950 (
            .O(N__35233),
            .I(N__35168));
    CascadeMux I__6949 (
            .O(N__35232),
            .I(N__35165));
    InMux I__6948 (
            .O(N__35231),
            .I(N__35150));
    InMux I__6947 (
            .O(N__35230),
            .I(N__35150));
    InMux I__6946 (
            .O(N__35229),
            .I(N__35150));
    InMux I__6945 (
            .O(N__35228),
            .I(N__35150));
    InMux I__6944 (
            .O(N__35227),
            .I(N__35150));
    InMux I__6943 (
            .O(N__35226),
            .I(N__35150));
    CascadeMux I__6942 (
            .O(N__35225),
            .I(N__35128));
    CascadeMux I__6941 (
            .O(N__35224),
            .I(N__35124));
    CascadeMux I__6940 (
            .O(N__35223),
            .I(N__35120));
    CascadeMux I__6939 (
            .O(N__35222),
            .I(N__35116));
    InMux I__6938 (
            .O(N__35221),
            .I(N__35093));
    InMux I__6937 (
            .O(N__35220),
            .I(N__35093));
    InMux I__6936 (
            .O(N__35219),
            .I(N__35093));
    InMux I__6935 (
            .O(N__35218),
            .I(N__35093));
    InMux I__6934 (
            .O(N__35217),
            .I(N__35093));
    InMux I__6933 (
            .O(N__35216),
            .I(N__35093));
    InMux I__6932 (
            .O(N__35215),
            .I(N__35093));
    LocalMux I__6931 (
            .O(N__35210),
            .I(N__35088));
    LocalMux I__6930 (
            .O(N__35199),
            .I(N__35088));
    InMux I__6929 (
            .O(N__35198),
            .I(N__35085));
    InMux I__6928 (
            .O(N__35197),
            .I(N__35080));
    InMux I__6927 (
            .O(N__35194),
            .I(N__35080));
    CascadeMux I__6926 (
            .O(N__35193),
            .I(N__35077));
    CascadeMux I__6925 (
            .O(N__35192),
            .I(N__35073));
    InMux I__6924 (
            .O(N__35189),
            .I(N__35069));
    InMux I__6923 (
            .O(N__35188),
            .I(N__35062));
    InMux I__6922 (
            .O(N__35187),
            .I(N__35062));
    InMux I__6921 (
            .O(N__35186),
            .I(N__35062));
    InMux I__6920 (
            .O(N__35185),
            .I(N__35057));
    InMux I__6919 (
            .O(N__35184),
            .I(N__35057));
    LocalMux I__6918 (
            .O(N__35181),
            .I(N__35054));
    InMux I__6917 (
            .O(N__35178),
            .I(N__35051));
    InMux I__6916 (
            .O(N__35177),
            .I(N__35038));
    InMux I__6915 (
            .O(N__35176),
            .I(N__35038));
    InMux I__6914 (
            .O(N__35175),
            .I(N__35038));
    InMux I__6913 (
            .O(N__35172),
            .I(N__35038));
    InMux I__6912 (
            .O(N__35171),
            .I(N__35038));
    InMux I__6911 (
            .O(N__35168),
            .I(N__35038));
    InMux I__6910 (
            .O(N__35165),
            .I(N__35031));
    InMux I__6909 (
            .O(N__35164),
            .I(N__35031));
    InMux I__6908 (
            .O(N__35163),
            .I(N__35031));
    LocalMux I__6907 (
            .O(N__35150),
            .I(N__35028));
    InMux I__6906 (
            .O(N__35149),
            .I(N__35023));
    InMux I__6905 (
            .O(N__35148),
            .I(N__35023));
    CascadeMux I__6904 (
            .O(N__35147),
            .I(N__35020));
    CascadeMux I__6903 (
            .O(N__35146),
            .I(N__35017));
    CascadeMux I__6902 (
            .O(N__35145),
            .I(N__35009));
    CascadeMux I__6901 (
            .O(N__35144),
            .I(N__35005));
    CascadeMux I__6900 (
            .O(N__35143),
            .I(N__35001));
    InMux I__6899 (
            .O(N__35142),
            .I(N__34993));
    InMux I__6898 (
            .O(N__35141),
            .I(N__34993));
    InMux I__6897 (
            .O(N__35140),
            .I(N__34993));
    CascadeMux I__6896 (
            .O(N__35139),
            .I(N__34990));
    CascadeMux I__6895 (
            .O(N__35138),
            .I(N__34986));
    CascadeMux I__6894 (
            .O(N__35137),
            .I(N__34982));
    CascadeMux I__6893 (
            .O(N__35136),
            .I(N__34978));
    InMux I__6892 (
            .O(N__35135),
            .I(N__34966));
    InMux I__6891 (
            .O(N__35134),
            .I(N__34966));
    InMux I__6890 (
            .O(N__35133),
            .I(N__34966));
    InMux I__6889 (
            .O(N__35132),
            .I(N__34966));
    InMux I__6888 (
            .O(N__35131),
            .I(N__34966));
    InMux I__6887 (
            .O(N__35128),
            .I(N__34949));
    InMux I__6886 (
            .O(N__35127),
            .I(N__34949));
    InMux I__6885 (
            .O(N__35124),
            .I(N__34949));
    InMux I__6884 (
            .O(N__35123),
            .I(N__34949));
    InMux I__6883 (
            .O(N__35120),
            .I(N__34949));
    InMux I__6882 (
            .O(N__35119),
            .I(N__34949));
    InMux I__6881 (
            .O(N__35116),
            .I(N__34949));
    InMux I__6880 (
            .O(N__35115),
            .I(N__34949));
    CascadeMux I__6879 (
            .O(N__35114),
            .I(N__34946));
    CascadeMux I__6878 (
            .O(N__35113),
            .I(N__34942));
    CascadeMux I__6877 (
            .O(N__35112),
            .I(N__34938));
    CascadeMux I__6876 (
            .O(N__35111),
            .I(N__34934));
    CascadeMux I__6875 (
            .O(N__35110),
            .I(N__34930));
    CascadeMux I__6874 (
            .O(N__35109),
            .I(N__34926));
    CascadeMux I__6873 (
            .O(N__35108),
            .I(N__34922));
    LocalMux I__6872 (
            .O(N__35093),
            .I(N__34918));
    Span4Mux_h I__6871 (
            .O(N__35088),
            .I(N__34911));
    LocalMux I__6870 (
            .O(N__35085),
            .I(N__34911));
    LocalMux I__6869 (
            .O(N__35080),
            .I(N__34911));
    InMux I__6868 (
            .O(N__35077),
            .I(N__34908));
    InMux I__6867 (
            .O(N__35076),
            .I(N__34903));
    InMux I__6866 (
            .O(N__35073),
            .I(N__34903));
    CascadeMux I__6865 (
            .O(N__35072),
            .I(N__34897));
    LocalMux I__6864 (
            .O(N__35069),
            .I(N__34890));
    LocalMux I__6863 (
            .O(N__35062),
            .I(N__34885));
    LocalMux I__6862 (
            .O(N__35057),
            .I(N__34885));
    Span4Mux_v I__6861 (
            .O(N__35054),
            .I(N__34876));
    LocalMux I__6860 (
            .O(N__35051),
            .I(N__34876));
    LocalMux I__6859 (
            .O(N__35038),
            .I(N__34876));
    LocalMux I__6858 (
            .O(N__35031),
            .I(N__34876));
    Span4Mux_h I__6857 (
            .O(N__35028),
            .I(N__34864));
    LocalMux I__6856 (
            .O(N__35023),
            .I(N__34864));
    InMux I__6855 (
            .O(N__35020),
            .I(N__34851));
    InMux I__6854 (
            .O(N__35017),
            .I(N__34851));
    InMux I__6853 (
            .O(N__35016),
            .I(N__34851));
    InMux I__6852 (
            .O(N__35015),
            .I(N__34851));
    InMux I__6851 (
            .O(N__35014),
            .I(N__34851));
    InMux I__6850 (
            .O(N__35013),
            .I(N__34851));
    InMux I__6849 (
            .O(N__35012),
            .I(N__34836));
    InMux I__6848 (
            .O(N__35009),
            .I(N__34836));
    InMux I__6847 (
            .O(N__35008),
            .I(N__34836));
    InMux I__6846 (
            .O(N__35005),
            .I(N__34836));
    InMux I__6845 (
            .O(N__35004),
            .I(N__34836));
    InMux I__6844 (
            .O(N__35001),
            .I(N__34836));
    InMux I__6843 (
            .O(N__35000),
            .I(N__34836));
    LocalMux I__6842 (
            .O(N__34993),
            .I(N__34833));
    InMux I__6841 (
            .O(N__34990),
            .I(N__34816));
    InMux I__6840 (
            .O(N__34989),
            .I(N__34816));
    InMux I__6839 (
            .O(N__34986),
            .I(N__34816));
    InMux I__6838 (
            .O(N__34985),
            .I(N__34816));
    InMux I__6837 (
            .O(N__34982),
            .I(N__34816));
    InMux I__6836 (
            .O(N__34981),
            .I(N__34816));
    InMux I__6835 (
            .O(N__34978),
            .I(N__34816));
    InMux I__6834 (
            .O(N__34977),
            .I(N__34816));
    LocalMux I__6833 (
            .O(N__34966),
            .I(N__34811));
    LocalMux I__6832 (
            .O(N__34949),
            .I(N__34811));
    InMux I__6831 (
            .O(N__34946),
            .I(N__34794));
    InMux I__6830 (
            .O(N__34945),
            .I(N__34794));
    InMux I__6829 (
            .O(N__34942),
            .I(N__34794));
    InMux I__6828 (
            .O(N__34941),
            .I(N__34794));
    InMux I__6827 (
            .O(N__34938),
            .I(N__34794));
    InMux I__6826 (
            .O(N__34937),
            .I(N__34794));
    InMux I__6825 (
            .O(N__34934),
            .I(N__34794));
    InMux I__6824 (
            .O(N__34933),
            .I(N__34794));
    InMux I__6823 (
            .O(N__34930),
            .I(N__34781));
    InMux I__6822 (
            .O(N__34929),
            .I(N__34781));
    InMux I__6821 (
            .O(N__34926),
            .I(N__34781));
    InMux I__6820 (
            .O(N__34925),
            .I(N__34781));
    InMux I__6819 (
            .O(N__34922),
            .I(N__34781));
    InMux I__6818 (
            .O(N__34921),
            .I(N__34781));
    Span4Mux_h I__6817 (
            .O(N__34918),
            .I(N__34772));
    Span4Mux_v I__6816 (
            .O(N__34911),
            .I(N__34772));
    LocalMux I__6815 (
            .O(N__34908),
            .I(N__34772));
    LocalMux I__6814 (
            .O(N__34903),
            .I(N__34772));
    InMux I__6813 (
            .O(N__34902),
            .I(N__34755));
    InMux I__6812 (
            .O(N__34901),
            .I(N__34755));
    InMux I__6811 (
            .O(N__34900),
            .I(N__34755));
    InMux I__6810 (
            .O(N__34897),
            .I(N__34755));
    InMux I__6809 (
            .O(N__34896),
            .I(N__34755));
    InMux I__6808 (
            .O(N__34895),
            .I(N__34755));
    InMux I__6807 (
            .O(N__34894),
            .I(N__34755));
    InMux I__6806 (
            .O(N__34893),
            .I(N__34755));
    Span4Mux_h I__6805 (
            .O(N__34890),
            .I(N__34750));
    Span4Mux_h I__6804 (
            .O(N__34885),
            .I(N__34750));
    Span4Mux_v I__6803 (
            .O(N__34876),
            .I(N__34747));
    CascadeMux I__6802 (
            .O(N__34875),
            .I(N__34744));
    CascadeMux I__6801 (
            .O(N__34874),
            .I(N__34740));
    CascadeMux I__6800 (
            .O(N__34873),
            .I(N__34736));
    CascadeMux I__6799 (
            .O(N__34872),
            .I(N__34732));
    CascadeMux I__6798 (
            .O(N__34871),
            .I(N__34728));
    CascadeMux I__6797 (
            .O(N__34870),
            .I(N__34724));
    CascadeMux I__6796 (
            .O(N__34869),
            .I(N__34720));
    Span4Mux_h I__6795 (
            .O(N__34864),
            .I(N__34702));
    LocalMux I__6794 (
            .O(N__34851),
            .I(N__34702));
    LocalMux I__6793 (
            .O(N__34836),
            .I(N__34702));
    Span4Mux_v I__6792 (
            .O(N__34833),
            .I(N__34702));
    LocalMux I__6791 (
            .O(N__34816),
            .I(N__34702));
    Span4Mux_v I__6790 (
            .O(N__34811),
            .I(N__34702));
    LocalMux I__6789 (
            .O(N__34794),
            .I(N__34702));
    LocalMux I__6788 (
            .O(N__34781),
            .I(N__34702));
    Span4Mux_v I__6787 (
            .O(N__34772),
            .I(N__34699));
    LocalMux I__6786 (
            .O(N__34755),
            .I(N__34696));
    Span4Mux_v I__6785 (
            .O(N__34750),
            .I(N__34691));
    Span4Mux_v I__6784 (
            .O(N__34747),
            .I(N__34691));
    InMux I__6783 (
            .O(N__34744),
            .I(N__34674));
    InMux I__6782 (
            .O(N__34743),
            .I(N__34674));
    InMux I__6781 (
            .O(N__34740),
            .I(N__34674));
    InMux I__6780 (
            .O(N__34739),
            .I(N__34674));
    InMux I__6779 (
            .O(N__34736),
            .I(N__34674));
    InMux I__6778 (
            .O(N__34735),
            .I(N__34674));
    InMux I__6777 (
            .O(N__34732),
            .I(N__34674));
    InMux I__6776 (
            .O(N__34731),
            .I(N__34674));
    InMux I__6775 (
            .O(N__34728),
            .I(N__34661));
    InMux I__6774 (
            .O(N__34727),
            .I(N__34661));
    InMux I__6773 (
            .O(N__34724),
            .I(N__34661));
    InMux I__6772 (
            .O(N__34723),
            .I(N__34661));
    InMux I__6771 (
            .O(N__34720),
            .I(N__34661));
    InMux I__6770 (
            .O(N__34719),
            .I(N__34661));
    Span4Mux_v I__6769 (
            .O(N__34702),
            .I(N__34658));
    Odrv4 I__6768 (
            .O(N__34699),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6767 (
            .O(N__34696),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6766 (
            .O(N__34691),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6765 (
            .O(N__34674),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6764 (
            .O(N__34661),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6763 (
            .O(N__34658),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__6762 (
            .O(N__34645),
            .I(N__34642));
    LocalMux I__6761 (
            .O(N__34642),
            .I(N__34639));
    Span4Mux_v I__6760 (
            .O(N__34639),
            .I(N__34634));
    InMux I__6759 (
            .O(N__34638),
            .I(N__34631));
    InMux I__6758 (
            .O(N__34637),
            .I(N__34628));
    Span4Mux_v I__6757 (
            .O(N__34634),
            .I(N__34623));
    LocalMux I__6756 (
            .O(N__34631),
            .I(N__34623));
    LocalMux I__6755 (
            .O(N__34628),
            .I(N__34620));
    Span4Mux_h I__6754 (
            .O(N__34623),
            .I(N__34617));
    Span12Mux_s11_h I__6753 (
            .O(N__34620),
            .I(N__34614));
    Odrv4 I__6752 (
            .O(N__34617),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv12 I__6751 (
            .O(N__34614),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__6750 (
            .O(N__34609),
            .I(N__34606));
    LocalMux I__6749 (
            .O(N__34606),
            .I(N__34603));
    Span4Mux_h I__6748 (
            .O(N__34603),
            .I(N__34600));
    Odrv4 I__6747 (
            .O(N__34600),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__6746 (
            .O(N__34597),
            .I(N__34594));
    LocalMux I__6745 (
            .O(N__34594),
            .I(N__34589));
    InMux I__6744 (
            .O(N__34593),
            .I(N__34586));
    InMux I__6743 (
            .O(N__34592),
            .I(N__34583));
    Span4Mux_v I__6742 (
            .O(N__34589),
            .I(N__34580));
    LocalMux I__6741 (
            .O(N__34586),
            .I(N__34577));
    LocalMux I__6740 (
            .O(N__34583),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__6739 (
            .O(N__34580),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__6738 (
            .O(N__34577),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__6737 (
            .O(N__34570),
            .I(N__34567));
    LocalMux I__6736 (
            .O(N__34567),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__6735 (
            .O(N__34564),
            .I(N__34560));
    InMux I__6734 (
            .O(N__34563),
            .I(N__34557));
    LocalMux I__6733 (
            .O(N__34560),
            .I(N__34551));
    LocalMux I__6732 (
            .O(N__34557),
            .I(N__34551));
    InMux I__6731 (
            .O(N__34556),
            .I(N__34548));
    Span4Mux_h I__6730 (
            .O(N__34551),
            .I(N__34545));
    LocalMux I__6729 (
            .O(N__34548),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__6728 (
            .O(N__34545),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__6727 (
            .O(N__34540),
            .I(N__34537));
    InMux I__6726 (
            .O(N__34537),
            .I(N__34534));
    LocalMux I__6725 (
            .O(N__34534),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__6724 (
            .O(N__34531),
            .I(N__34528));
    LocalMux I__6723 (
            .O(N__34528),
            .I(N__34523));
    InMux I__6722 (
            .O(N__34527),
            .I(N__34520));
    InMux I__6721 (
            .O(N__34526),
            .I(N__34517));
    Span4Mux_v I__6720 (
            .O(N__34523),
            .I(N__34514));
    LocalMux I__6719 (
            .O(N__34520),
            .I(N__34511));
    LocalMux I__6718 (
            .O(N__34517),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__6717 (
            .O(N__34514),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__6716 (
            .O(N__34511),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    CascadeMux I__6715 (
            .O(N__34504),
            .I(N__34501));
    InMux I__6714 (
            .O(N__34501),
            .I(N__34498));
    LocalMux I__6713 (
            .O(N__34498),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__6712 (
            .O(N__34495),
            .I(N__34490));
    InMux I__6711 (
            .O(N__34494),
            .I(N__34487));
    InMux I__6710 (
            .O(N__34493),
            .I(N__34484));
    LocalMux I__6709 (
            .O(N__34490),
            .I(N__34479));
    LocalMux I__6708 (
            .O(N__34487),
            .I(N__34479));
    LocalMux I__6707 (
            .O(N__34484),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__6706 (
            .O(N__34479),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__6705 (
            .O(N__34474),
            .I(N__34471));
    LocalMux I__6704 (
            .O(N__34471),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__6703 (
            .O(N__34468),
            .I(N__34463));
    InMux I__6702 (
            .O(N__34467),
            .I(N__34460));
    InMux I__6701 (
            .O(N__34466),
            .I(N__34457));
    LocalMux I__6700 (
            .O(N__34463),
            .I(N__34452));
    LocalMux I__6699 (
            .O(N__34460),
            .I(N__34452));
    LocalMux I__6698 (
            .O(N__34457),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__6697 (
            .O(N__34452),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    CascadeMux I__6696 (
            .O(N__34447),
            .I(N__34444));
    InMux I__6695 (
            .O(N__34444),
            .I(N__34441));
    LocalMux I__6694 (
            .O(N__34441),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__6693 (
            .O(N__34438),
            .I(N__34433));
    InMux I__6692 (
            .O(N__34437),
            .I(N__34430));
    InMux I__6691 (
            .O(N__34436),
            .I(N__34427));
    LocalMux I__6690 (
            .O(N__34433),
            .I(N__34424));
    LocalMux I__6689 (
            .O(N__34430),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__6688 (
            .O(N__34427),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__6687 (
            .O(N__34424),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__6686 (
            .O(N__34417),
            .I(N__34414));
    LocalMux I__6685 (
            .O(N__34414),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__6684 (
            .O(N__34411),
            .I(N__34408));
    LocalMux I__6683 (
            .O(N__34408),
            .I(N__34404));
    InMux I__6682 (
            .O(N__34407),
            .I(N__34401));
    Span4Mux_h I__6681 (
            .O(N__34404),
            .I(N__34398));
    LocalMux I__6680 (
            .O(N__34401),
            .I(N__34395));
    Span4Mux_h I__6679 (
            .O(N__34398),
            .I(N__34392));
    Span12Mux_s7_h I__6678 (
            .O(N__34395),
            .I(N__34389));
    Odrv4 I__6677 (
            .O(N__34392),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv12 I__6676 (
            .O(N__34389),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6675 (
            .O(N__34384),
            .I(N__34380));
    InMux I__6674 (
            .O(N__34383),
            .I(N__34377));
    LocalMux I__6673 (
            .O(N__34380),
            .I(N__34374));
    LocalMux I__6672 (
            .O(N__34377),
            .I(N__34371));
    Span4Mux_h I__6671 (
            .O(N__34374),
            .I(N__34368));
    Span4Mux_s3_h I__6670 (
            .O(N__34371),
            .I(N__34365));
    Span4Mux_h I__6669 (
            .O(N__34368),
            .I(N__34362));
    Span4Mux_h I__6668 (
            .O(N__34365),
            .I(N__34359));
    Odrv4 I__6667 (
            .O(N__34362),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__6666 (
            .O(N__34359),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__6665 (
            .O(N__34354),
            .I(N__34350));
    InMux I__6664 (
            .O(N__34353),
            .I(N__34347));
    LocalMux I__6663 (
            .O(N__34350),
            .I(N__34344));
    LocalMux I__6662 (
            .O(N__34347),
            .I(N__34341));
    Sp12to4 I__6661 (
            .O(N__34344),
            .I(N__34338));
    Span12Mux_v I__6660 (
            .O(N__34341),
            .I(N__34333));
    Span12Mux_v I__6659 (
            .O(N__34338),
            .I(N__34333));
    Odrv12 I__6658 (
            .O(N__34333),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__6657 (
            .O(N__34330),
            .I(N__34326));
    InMux I__6656 (
            .O(N__34329),
            .I(N__34323));
    LocalMux I__6655 (
            .O(N__34326),
            .I(N__34320));
    LocalMux I__6654 (
            .O(N__34323),
            .I(N__34317));
    Span4Mux_s3_h I__6653 (
            .O(N__34320),
            .I(N__34314));
    Span4Mux_v I__6652 (
            .O(N__34317),
            .I(N__34311));
    Sp12to4 I__6651 (
            .O(N__34314),
            .I(N__34308));
    Sp12to4 I__6650 (
            .O(N__34311),
            .I(N__34303));
    Span12Mux_v I__6649 (
            .O(N__34308),
            .I(N__34303));
    Odrv12 I__6648 (
            .O(N__34303),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__6647 (
            .O(N__34300),
            .I(N__34296));
    InMux I__6646 (
            .O(N__34299),
            .I(N__34293));
    LocalMux I__6645 (
            .O(N__34296),
            .I(N__34290));
    LocalMux I__6644 (
            .O(N__34293),
            .I(N__34287));
    Span4Mux_v I__6643 (
            .O(N__34290),
            .I(N__34284));
    Span4Mux_v I__6642 (
            .O(N__34287),
            .I(N__34281));
    Span4Mux_h I__6641 (
            .O(N__34284),
            .I(N__34276));
    Span4Mux_h I__6640 (
            .O(N__34281),
            .I(N__34276));
    Odrv4 I__6639 (
            .O(N__34276),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__6638 (
            .O(N__34273),
            .I(N__34269));
    InMux I__6637 (
            .O(N__34272),
            .I(N__34266));
    LocalMux I__6636 (
            .O(N__34269),
            .I(N__34263));
    LocalMux I__6635 (
            .O(N__34266),
            .I(N__34260));
    Span4Mux_s2_h I__6634 (
            .O(N__34263),
            .I(N__34257));
    Span4Mux_v I__6633 (
            .O(N__34260),
            .I(N__34254));
    Sp12to4 I__6632 (
            .O(N__34257),
            .I(N__34251));
    Sp12to4 I__6631 (
            .O(N__34254),
            .I(N__34246));
    Span12Mux_v I__6630 (
            .O(N__34251),
            .I(N__34246));
    Odrv12 I__6629 (
            .O(N__34246),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__6628 (
            .O(N__34243),
            .I(N__34239));
    InMux I__6627 (
            .O(N__34242),
            .I(N__34236));
    LocalMux I__6626 (
            .O(N__34239),
            .I(N__34233));
    LocalMux I__6625 (
            .O(N__34236),
            .I(N__34230));
    Span4Mux_v I__6624 (
            .O(N__34233),
            .I(N__34227));
    Span4Mux_h I__6623 (
            .O(N__34230),
            .I(N__34224));
    Sp12to4 I__6622 (
            .O(N__34227),
            .I(N__34221));
    Span4Mux_h I__6621 (
            .O(N__34224),
            .I(N__34218));
    Span12Mux_s7_h I__6620 (
            .O(N__34221),
            .I(N__34215));
    Odrv4 I__6619 (
            .O(N__34218),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv12 I__6618 (
            .O(N__34215),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__6617 (
            .O(N__34210),
            .I(N__34206));
    InMux I__6616 (
            .O(N__34209),
            .I(N__34203));
    LocalMux I__6615 (
            .O(N__34206),
            .I(N__34200));
    LocalMux I__6614 (
            .O(N__34203),
            .I(N__34197));
    Span4Mux_v I__6613 (
            .O(N__34200),
            .I(N__34194));
    Span4Mux_h I__6612 (
            .O(N__34197),
            .I(N__34191));
    Sp12to4 I__6611 (
            .O(N__34194),
            .I(N__34188));
    Span4Mux_h I__6610 (
            .O(N__34191),
            .I(N__34185));
    Span12Mux_s7_h I__6609 (
            .O(N__34188),
            .I(N__34182));
    Odrv4 I__6608 (
            .O(N__34185),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv12 I__6607 (
            .O(N__34182),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__6606 (
            .O(N__34177),
            .I(N__34173));
    InMux I__6605 (
            .O(N__34176),
            .I(N__34170));
    LocalMux I__6604 (
            .O(N__34173),
            .I(N__34167));
    LocalMux I__6603 (
            .O(N__34170),
            .I(N__34164));
    Span4Mux_v I__6602 (
            .O(N__34167),
            .I(N__34161));
    Span4Mux_h I__6601 (
            .O(N__34164),
            .I(N__34158));
    Sp12to4 I__6600 (
            .O(N__34161),
            .I(N__34155));
    Span4Mux_h I__6599 (
            .O(N__34158),
            .I(N__34152));
    Span12Mux_s7_h I__6598 (
            .O(N__34155),
            .I(N__34149));
    Odrv4 I__6597 (
            .O(N__34152),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv12 I__6596 (
            .O(N__34149),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    IoInMux I__6595 (
            .O(N__34144),
            .I(N__34141));
    LocalMux I__6594 (
            .O(N__34141),
            .I(N__34138));
    Span12Mux_s10_v I__6593 (
            .O(N__34138),
            .I(N__34135));
    Odrv12 I__6592 (
            .O(N__34135),
            .I(s2_phy_c));
    InMux I__6591 (
            .O(N__34132),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__6590 (
            .O(N__34129),
            .I(N__34124));
    InMux I__6589 (
            .O(N__34128),
            .I(N__34121));
    InMux I__6588 (
            .O(N__34127),
            .I(N__34118));
    LocalMux I__6587 (
            .O(N__34124),
            .I(N__34115));
    LocalMux I__6586 (
            .O(N__34121),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__6585 (
            .O(N__34118),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__6584 (
            .O(N__34115),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__6583 (
            .O(N__34108),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__6582 (
            .O(N__34105),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__6581 (
            .O(N__34102),
            .I(N__34099));
    InMux I__6580 (
            .O(N__34099),
            .I(N__34094));
    InMux I__6579 (
            .O(N__34098),
            .I(N__34091));
    InMux I__6578 (
            .O(N__34097),
            .I(N__34088));
    LocalMux I__6577 (
            .O(N__34094),
            .I(N__34085));
    LocalMux I__6576 (
            .O(N__34091),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__6575 (
            .O(N__34088),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv12 I__6574 (
            .O(N__34085),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__6573 (
            .O(N__34078),
            .I(N__34074));
    InMux I__6572 (
            .O(N__34077),
            .I(N__34071));
    LocalMux I__6571 (
            .O(N__34074),
            .I(N__34068));
    LocalMux I__6570 (
            .O(N__34071),
            .I(N__34065));
    Span4Mux_h I__6569 (
            .O(N__34068),
            .I(N__34062));
    Span4Mux_v I__6568 (
            .O(N__34065),
            .I(N__34059));
    Span4Mux_h I__6567 (
            .O(N__34062),
            .I(N__34056));
    Sp12to4 I__6566 (
            .O(N__34059),
            .I(N__34053));
    Odrv4 I__6565 (
            .O(N__34056),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__6564 (
            .O(N__34053),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__6563 (
            .O(N__34048),
            .I(N__34044));
    InMux I__6562 (
            .O(N__34047),
            .I(N__34041));
    LocalMux I__6561 (
            .O(N__34044),
            .I(N__34038));
    LocalMux I__6560 (
            .O(N__34041),
            .I(N__34035));
    Span4Mux_h I__6559 (
            .O(N__34038),
            .I(N__34032));
    Span4Mux_s3_h I__6558 (
            .O(N__34035),
            .I(N__34029));
    Span4Mux_h I__6557 (
            .O(N__34032),
            .I(N__34024));
    Span4Mux_h I__6556 (
            .O(N__34029),
            .I(N__34024));
    Odrv4 I__6555 (
            .O(N__34024),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__6554 (
            .O(N__34021),
            .I(N__34018));
    LocalMux I__6553 (
            .O(N__34018),
            .I(N__34015));
    Span4Mux_v I__6552 (
            .O(N__34015),
            .I(N__34011));
    InMux I__6551 (
            .O(N__34014),
            .I(N__34008));
    Sp12to4 I__6550 (
            .O(N__34011),
            .I(N__34005));
    LocalMux I__6549 (
            .O(N__34008),
            .I(N__34002));
    Span12Mux_s7_h I__6548 (
            .O(N__34005),
            .I(N__33999));
    Odrv12 I__6547 (
            .O(N__34002),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__6546 (
            .O(N__33999),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__6545 (
            .O(N__33994),
            .I(N__33990));
    InMux I__6544 (
            .O(N__33993),
            .I(N__33987));
    LocalMux I__6543 (
            .O(N__33990),
            .I(N__33984));
    LocalMux I__6542 (
            .O(N__33987),
            .I(N__33981));
    Span4Mux_v I__6541 (
            .O(N__33984),
            .I(N__33978));
    Span4Mux_v I__6540 (
            .O(N__33981),
            .I(N__33975));
    Span4Mux_h I__6539 (
            .O(N__33978),
            .I(N__33972));
    Span4Mux_h I__6538 (
            .O(N__33975),
            .I(N__33969));
    Odrv4 I__6537 (
            .O(N__33972),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__6536 (
            .O(N__33969),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__6535 (
            .O(N__33964),
            .I(N__33961));
    LocalMux I__6534 (
            .O(N__33961),
            .I(N__33957));
    InMux I__6533 (
            .O(N__33960),
            .I(N__33954));
    Span4Mux_h I__6532 (
            .O(N__33957),
            .I(N__33951));
    LocalMux I__6531 (
            .O(N__33954),
            .I(N__33948));
    Span4Mux_h I__6530 (
            .O(N__33951),
            .I(N__33945));
    Span12Mux_s7_h I__6529 (
            .O(N__33948),
            .I(N__33942));
    Odrv4 I__6528 (
            .O(N__33945),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    Odrv12 I__6527 (
            .O(N__33942),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__6526 (
            .O(N__33937),
            .I(N__33933));
    InMux I__6525 (
            .O(N__33936),
            .I(N__33930));
    LocalMux I__6524 (
            .O(N__33933),
            .I(N__33927));
    LocalMux I__6523 (
            .O(N__33930),
            .I(N__33924));
    Span4Mux_v I__6522 (
            .O(N__33927),
            .I(N__33921));
    Span4Mux_v I__6521 (
            .O(N__33924),
            .I(N__33918));
    Sp12to4 I__6520 (
            .O(N__33921),
            .I(N__33915));
    Span4Mux_h I__6519 (
            .O(N__33918),
            .I(N__33912));
    Span12Mux_s7_h I__6518 (
            .O(N__33915),
            .I(N__33909));
    Odrv4 I__6517 (
            .O(N__33912),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv12 I__6516 (
            .O(N__33909),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    CascadeMux I__6515 (
            .O(N__33904),
            .I(N__33900));
    InMux I__6514 (
            .O(N__33903),
            .I(N__33895));
    InMux I__6513 (
            .O(N__33900),
            .I(N__33895));
    LocalMux I__6512 (
            .O(N__33895),
            .I(N__33891));
    InMux I__6511 (
            .O(N__33894),
            .I(N__33888));
    Span4Mux_v I__6510 (
            .O(N__33891),
            .I(N__33885));
    LocalMux I__6509 (
            .O(N__33888),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__6508 (
            .O(N__33885),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__6507 (
            .O(N__33880),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__6506 (
            .O(N__33877),
            .I(N__33874));
    InMux I__6505 (
            .O(N__33874),
            .I(N__33867));
    InMux I__6504 (
            .O(N__33873),
            .I(N__33867));
    InMux I__6503 (
            .O(N__33872),
            .I(N__33864));
    LocalMux I__6502 (
            .O(N__33867),
            .I(N__33861));
    LocalMux I__6501 (
            .O(N__33864),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__6500 (
            .O(N__33861),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__6499 (
            .O(N__33856),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__6498 (
            .O(N__33853),
            .I(N__33846));
    InMux I__6497 (
            .O(N__33852),
            .I(N__33846));
    InMux I__6496 (
            .O(N__33851),
            .I(N__33843));
    LocalMux I__6495 (
            .O(N__33846),
            .I(N__33840));
    LocalMux I__6494 (
            .O(N__33843),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__6493 (
            .O(N__33840),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__6492 (
            .O(N__33835),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    CascadeMux I__6491 (
            .O(N__33832),
            .I(N__33829));
    InMux I__6490 (
            .O(N__33829),
            .I(N__33823));
    InMux I__6489 (
            .O(N__33828),
            .I(N__33823));
    LocalMux I__6488 (
            .O(N__33823),
            .I(N__33819));
    InMux I__6487 (
            .O(N__33822),
            .I(N__33816));
    Span4Mux_h I__6486 (
            .O(N__33819),
            .I(N__33813));
    LocalMux I__6485 (
            .O(N__33816),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__6484 (
            .O(N__33813),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__6483 (
            .O(N__33808),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__6482 (
            .O(N__33805),
            .I(N__33798));
    InMux I__6481 (
            .O(N__33804),
            .I(N__33798));
    InMux I__6480 (
            .O(N__33803),
            .I(N__33795));
    LocalMux I__6479 (
            .O(N__33798),
            .I(N__33792));
    LocalMux I__6478 (
            .O(N__33795),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__6477 (
            .O(N__33792),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__6476 (
            .O(N__33787),
            .I(bfn_13_15_0_));
    InMux I__6475 (
            .O(N__33784),
            .I(N__33779));
    InMux I__6474 (
            .O(N__33783),
            .I(N__33774));
    InMux I__6473 (
            .O(N__33782),
            .I(N__33774));
    LocalMux I__6472 (
            .O(N__33779),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__6471 (
            .O(N__33774),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__6470 (
            .O(N__33769),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    CascadeMux I__6469 (
            .O(N__33766),
            .I(N__33762));
    InMux I__6468 (
            .O(N__33765),
            .I(N__33758));
    InMux I__6467 (
            .O(N__33762),
            .I(N__33753));
    InMux I__6466 (
            .O(N__33761),
            .I(N__33753));
    LocalMux I__6465 (
            .O(N__33758),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__6464 (
            .O(N__33753),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__6463 (
            .O(N__33748),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    CascadeMux I__6462 (
            .O(N__33745),
            .I(N__33740));
    InMux I__6461 (
            .O(N__33744),
            .I(N__33737));
    InMux I__6460 (
            .O(N__33743),
            .I(N__33732));
    InMux I__6459 (
            .O(N__33740),
            .I(N__33732));
    LocalMux I__6458 (
            .O(N__33737),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__6457 (
            .O(N__33732),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__6456 (
            .O(N__33727),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__6455 (
            .O(N__33724),
            .I(N__33719));
    InMux I__6454 (
            .O(N__33723),
            .I(N__33714));
    InMux I__6453 (
            .O(N__33722),
            .I(N__33714));
    LocalMux I__6452 (
            .O(N__33719),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__6451 (
            .O(N__33714),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__6450 (
            .O(N__33709),
            .I(N__33705));
    InMux I__6449 (
            .O(N__33708),
            .I(N__33702));
    LocalMux I__6448 (
            .O(N__33705),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__6447 (
            .O(N__33702),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__6446 (
            .O(N__33697),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__6445 (
            .O(N__33694),
            .I(N__33690));
    InMux I__6444 (
            .O(N__33693),
            .I(N__33687));
    LocalMux I__6443 (
            .O(N__33690),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__6442 (
            .O(N__33687),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__6441 (
            .O(N__33682),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__6440 (
            .O(N__33679),
            .I(N__33675));
    InMux I__6439 (
            .O(N__33678),
            .I(N__33672));
    LocalMux I__6438 (
            .O(N__33675),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__6437 (
            .O(N__33672),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__6436 (
            .O(N__33667),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__6435 (
            .O(N__33664),
            .I(N__33658));
    InMux I__6434 (
            .O(N__33663),
            .I(N__33658));
    LocalMux I__6433 (
            .O(N__33658),
            .I(N__33654));
    InMux I__6432 (
            .O(N__33657),
            .I(N__33651));
    Span4Mux_h I__6431 (
            .O(N__33654),
            .I(N__33648));
    LocalMux I__6430 (
            .O(N__33651),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__6429 (
            .O(N__33648),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__6428 (
            .O(N__33643),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    CascadeMux I__6427 (
            .O(N__33640),
            .I(N__33637));
    InMux I__6426 (
            .O(N__33637),
            .I(N__33631));
    InMux I__6425 (
            .O(N__33636),
            .I(N__33631));
    LocalMux I__6424 (
            .O(N__33631),
            .I(N__33627));
    InMux I__6423 (
            .O(N__33630),
            .I(N__33624));
    Span4Mux_h I__6422 (
            .O(N__33627),
            .I(N__33621));
    LocalMux I__6421 (
            .O(N__33624),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__6420 (
            .O(N__33621),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__6419 (
            .O(N__33616),
            .I(bfn_13_14_0_));
    CascadeMux I__6418 (
            .O(N__33613),
            .I(N__33610));
    InMux I__6417 (
            .O(N__33610),
            .I(N__33604));
    InMux I__6416 (
            .O(N__33609),
            .I(N__33604));
    LocalMux I__6415 (
            .O(N__33604),
            .I(N__33600));
    InMux I__6414 (
            .O(N__33603),
            .I(N__33597));
    Span4Mux_v I__6413 (
            .O(N__33600),
            .I(N__33594));
    LocalMux I__6412 (
            .O(N__33597),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__6411 (
            .O(N__33594),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__6410 (
            .O(N__33589),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__6409 (
            .O(N__33586),
            .I(N__33580));
    InMux I__6408 (
            .O(N__33585),
            .I(N__33580));
    LocalMux I__6407 (
            .O(N__33580),
            .I(N__33576));
    InMux I__6406 (
            .O(N__33579),
            .I(N__33573));
    Span4Mux_h I__6405 (
            .O(N__33576),
            .I(N__33570));
    LocalMux I__6404 (
            .O(N__33573),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__6403 (
            .O(N__33570),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__6402 (
            .O(N__33565),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__6401 (
            .O(N__33562),
            .I(N__33555));
    InMux I__6400 (
            .O(N__33561),
            .I(N__33555));
    InMux I__6399 (
            .O(N__33560),
            .I(N__33552));
    LocalMux I__6398 (
            .O(N__33555),
            .I(N__33549));
    LocalMux I__6397 (
            .O(N__33552),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__6396 (
            .O(N__33549),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__6395 (
            .O(N__33544),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__6394 (
            .O(N__33541),
            .I(N__33537));
    InMux I__6393 (
            .O(N__33540),
            .I(N__33534));
    LocalMux I__6392 (
            .O(N__33537),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__6391 (
            .O(N__33534),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__6390 (
            .O(N__33529),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__6389 (
            .O(N__33526),
            .I(N__33522));
    InMux I__6388 (
            .O(N__33525),
            .I(N__33519));
    LocalMux I__6387 (
            .O(N__33522),
            .I(N__33516));
    LocalMux I__6386 (
            .O(N__33519),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__6385 (
            .O(N__33516),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__6384 (
            .O(N__33511),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__6383 (
            .O(N__33508),
            .I(N__33504));
    InMux I__6382 (
            .O(N__33507),
            .I(N__33501));
    LocalMux I__6381 (
            .O(N__33504),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__6380 (
            .O(N__33501),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__6379 (
            .O(N__33496),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__6378 (
            .O(N__33493),
            .I(N__33489));
    InMux I__6377 (
            .O(N__33492),
            .I(N__33486));
    LocalMux I__6376 (
            .O(N__33489),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__6375 (
            .O(N__33486),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__6374 (
            .O(N__33481),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__6373 (
            .O(N__33478),
            .I(N__33474));
    InMux I__6372 (
            .O(N__33477),
            .I(N__33471));
    LocalMux I__6371 (
            .O(N__33474),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__6370 (
            .O(N__33471),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__6369 (
            .O(N__33466),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__6368 (
            .O(N__33463),
            .I(N__33459));
    InMux I__6367 (
            .O(N__33462),
            .I(N__33456));
    LocalMux I__6366 (
            .O(N__33459),
            .I(N__33453));
    LocalMux I__6365 (
            .O(N__33456),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__6364 (
            .O(N__33453),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__6363 (
            .O(N__33448),
            .I(bfn_13_13_0_));
    InMux I__6362 (
            .O(N__33445),
            .I(N__33441));
    InMux I__6361 (
            .O(N__33444),
            .I(N__33438));
    LocalMux I__6360 (
            .O(N__33441),
            .I(N__33435));
    LocalMux I__6359 (
            .O(N__33438),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__6358 (
            .O(N__33435),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__6357 (
            .O(N__33430),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__6356 (
            .O(N__33427),
            .I(N__33423));
    InMux I__6355 (
            .O(N__33426),
            .I(N__33420));
    LocalMux I__6354 (
            .O(N__33423),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__6353 (
            .O(N__33420),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__6352 (
            .O(N__33415),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__6351 (
            .O(N__33412),
            .I(N__33408));
    InMux I__6350 (
            .O(N__33411),
            .I(N__33405));
    LocalMux I__6349 (
            .O(N__33408),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__6348 (
            .O(N__33405),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__6347 (
            .O(N__33400),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__6346 (
            .O(N__33397),
            .I(N__33391));
    InMux I__6345 (
            .O(N__33396),
            .I(N__33391));
    LocalMux I__6344 (
            .O(N__33391),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__6343 (
            .O(N__33388),
            .I(N__33382));
    InMux I__6342 (
            .O(N__33387),
            .I(N__33382));
    LocalMux I__6341 (
            .O(N__33382),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__6340 (
            .O(N__33379),
            .I(N__33375));
    InMux I__6339 (
            .O(N__33378),
            .I(N__33372));
    LocalMux I__6338 (
            .O(N__33375),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__6337 (
            .O(N__33372),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__6336 (
            .O(N__33367),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__6335 (
            .O(N__33364),
            .I(N__33361));
    InMux I__6334 (
            .O(N__33361),
            .I(N__33357));
    InMux I__6333 (
            .O(N__33360),
            .I(N__33354));
    LocalMux I__6332 (
            .O(N__33357),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__6331 (
            .O(N__33354),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__6330 (
            .O(N__33349),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__6329 (
            .O(N__33346),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__6328 (
            .O(N__33343),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__6327 (
            .O(N__33340),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__6326 (
            .O(N__33337),
            .I(bfn_13_10_0_));
    InMux I__6325 (
            .O(N__33334),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__6324 (
            .O(N__33331),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__6323 (
            .O(N__33328),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__6322 (
            .O(N__33325),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6321 (
            .O(N__33322),
            .I(N__33284));
    InMux I__6320 (
            .O(N__33321),
            .I(N__33284));
    InMux I__6319 (
            .O(N__33320),
            .I(N__33284));
    InMux I__6318 (
            .O(N__33319),
            .I(N__33284));
    InMux I__6317 (
            .O(N__33318),
            .I(N__33275));
    InMux I__6316 (
            .O(N__33317),
            .I(N__33275));
    InMux I__6315 (
            .O(N__33316),
            .I(N__33275));
    InMux I__6314 (
            .O(N__33315),
            .I(N__33275));
    InMux I__6313 (
            .O(N__33314),
            .I(N__33268));
    InMux I__6312 (
            .O(N__33313),
            .I(N__33268));
    InMux I__6311 (
            .O(N__33312),
            .I(N__33268));
    InMux I__6310 (
            .O(N__33311),
            .I(N__33259));
    InMux I__6309 (
            .O(N__33310),
            .I(N__33259));
    InMux I__6308 (
            .O(N__33309),
            .I(N__33259));
    InMux I__6307 (
            .O(N__33308),
            .I(N__33259));
    InMux I__6306 (
            .O(N__33307),
            .I(N__33252));
    InMux I__6305 (
            .O(N__33306),
            .I(N__33252));
    InMux I__6304 (
            .O(N__33305),
            .I(N__33252));
    InMux I__6303 (
            .O(N__33304),
            .I(N__33243));
    InMux I__6302 (
            .O(N__33303),
            .I(N__33243));
    InMux I__6301 (
            .O(N__33302),
            .I(N__33243));
    InMux I__6300 (
            .O(N__33301),
            .I(N__33243));
    InMux I__6299 (
            .O(N__33300),
            .I(N__33234));
    InMux I__6298 (
            .O(N__33299),
            .I(N__33234));
    InMux I__6297 (
            .O(N__33298),
            .I(N__33234));
    InMux I__6296 (
            .O(N__33297),
            .I(N__33234));
    InMux I__6295 (
            .O(N__33296),
            .I(N__33225));
    InMux I__6294 (
            .O(N__33295),
            .I(N__33225));
    InMux I__6293 (
            .O(N__33294),
            .I(N__33225));
    InMux I__6292 (
            .O(N__33293),
            .I(N__33225));
    LocalMux I__6291 (
            .O(N__33284),
            .I(N__33220));
    LocalMux I__6290 (
            .O(N__33275),
            .I(N__33220));
    LocalMux I__6289 (
            .O(N__33268),
            .I(N__33215));
    LocalMux I__6288 (
            .O(N__33259),
            .I(N__33215));
    LocalMux I__6287 (
            .O(N__33252),
            .I(N__33208));
    LocalMux I__6286 (
            .O(N__33243),
            .I(N__33208));
    LocalMux I__6285 (
            .O(N__33234),
            .I(N__33208));
    LocalMux I__6284 (
            .O(N__33225),
            .I(N__33205));
    Span4Mux_h I__6283 (
            .O(N__33220),
            .I(N__33198));
    Span4Mux_v I__6282 (
            .O(N__33215),
            .I(N__33198));
    Span4Mux_v I__6281 (
            .O(N__33208),
            .I(N__33198));
    Span4Mux_h I__6280 (
            .O(N__33205),
            .I(N__33195));
    Odrv4 I__6279 (
            .O(N__33198),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6278 (
            .O(N__33195),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__6277 (
            .O(N__33190),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__6276 (
            .O(N__33187),
            .I(N__33183));
    CEMux I__6275 (
            .O(N__33186),
            .I(N__33178));
    LocalMux I__6274 (
            .O(N__33183),
            .I(N__33175));
    CEMux I__6273 (
            .O(N__33182),
            .I(N__33172));
    CEMux I__6272 (
            .O(N__33181),
            .I(N__33169));
    LocalMux I__6271 (
            .O(N__33178),
            .I(N__33166));
    Span4Mux_h I__6270 (
            .O(N__33175),
            .I(N__33163));
    LocalMux I__6269 (
            .O(N__33172),
            .I(N__33160));
    LocalMux I__6268 (
            .O(N__33169),
            .I(N__33157));
    Span4Mux_v I__6267 (
            .O(N__33166),
            .I(N__33154));
    Span4Mux_v I__6266 (
            .O(N__33163),
            .I(N__33151));
    Span4Mux_h I__6265 (
            .O(N__33160),
            .I(N__33148));
    Span4Mux_v I__6264 (
            .O(N__33157),
            .I(N__33143));
    Span4Mux_h I__6263 (
            .O(N__33154),
            .I(N__33143));
    Odrv4 I__6262 (
            .O(N__33151),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    Odrv4 I__6261 (
            .O(N__33148),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    Odrv4 I__6260 (
            .O(N__33143),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    InMux I__6259 (
            .O(N__33136),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__6258 (
            .O(N__33133),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__6257 (
            .O(N__33130),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__6256 (
            .O(N__33127),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__6255 (
            .O(N__33124),
            .I(bfn_13_9_0_));
    InMux I__6254 (
            .O(N__33121),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__6253 (
            .O(N__33118),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6252 (
            .O(N__33115),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__6251 (
            .O(N__33112),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__6250 (
            .O(N__33109),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__6249 (
            .O(N__33106),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__6248 (
            .O(N__33103),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__6247 (
            .O(N__33100),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__6246 (
            .O(N__33097),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__6245 (
            .O(N__33094),
            .I(bfn_13_8_0_));
    InMux I__6244 (
            .O(N__33091),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__6243 (
            .O(N__33088),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6242 (
            .O(N__33085),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__6241 (
            .O(N__33082),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__6240 (
            .O(N__33079),
            .I(bfn_12_27_0_));
    InMux I__6239 (
            .O(N__33076),
            .I(N__33062));
    InMux I__6238 (
            .O(N__33075),
            .I(N__33062));
    InMux I__6237 (
            .O(N__33074),
            .I(N__33053));
    InMux I__6236 (
            .O(N__33073),
            .I(N__33053));
    InMux I__6235 (
            .O(N__33072),
            .I(N__33053));
    InMux I__6234 (
            .O(N__33071),
            .I(N__33053));
    InMux I__6233 (
            .O(N__33070),
            .I(N__33044));
    InMux I__6232 (
            .O(N__33069),
            .I(N__33044));
    InMux I__6231 (
            .O(N__33068),
            .I(N__33044));
    InMux I__6230 (
            .O(N__33067),
            .I(N__33044));
    LocalMux I__6229 (
            .O(N__33062),
            .I(N__33041));
    LocalMux I__6228 (
            .O(N__33053),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__6227 (
            .O(N__33044),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__6226 (
            .O(N__33041),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__6225 (
            .O(N__33034),
            .I(\pwm_generator_inst.counter_cry_8 ));
    IoInMux I__6224 (
            .O(N__33031),
            .I(N__33028));
    LocalMux I__6223 (
            .O(N__33028),
            .I(N__33025));
    IoSpan4Mux I__6222 (
            .O(N__33025),
            .I(N__33022));
    Span4Mux_s0_v I__6221 (
            .O(N__33022),
            .I(N__33019));
    Odrv4 I__6220 (
            .O(N__33019),
            .I(GB_BUFFER_red_c_g_THRU_CO));
    InMux I__6219 (
            .O(N__33016),
            .I(bfn_13_7_0_));
    InMux I__6218 (
            .O(N__33013),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__6217 (
            .O(N__33010),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__6216 (
            .O(N__33007),
            .I(N__33004));
    LocalMux I__6215 (
            .O(N__33004),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    CascadeMux I__6214 (
            .O(N__33001),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__6213 (
            .O(N__32998),
            .I(bfn_12_26_0_));
    InMux I__6212 (
            .O(N__32995),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__6211 (
            .O(N__32992),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__6210 (
            .O(N__32989),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__6209 (
            .O(N__32986),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__6208 (
            .O(N__32983),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__6207 (
            .O(N__32980),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__6206 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__6205 (
            .O(N__32974),
            .I(N__32971));
    Span4Mux_h I__6204 (
            .O(N__32971),
            .I(N__32966));
    InMux I__6203 (
            .O(N__32970),
            .I(N__32963));
    InMux I__6202 (
            .O(N__32969),
            .I(N__32960));
    Odrv4 I__6201 (
            .O(N__32966),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__6200 (
            .O(N__32963),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__6199 (
            .O(N__32960),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__6198 (
            .O(N__32953),
            .I(N__32949));
    InMux I__6197 (
            .O(N__32952),
            .I(N__32946));
    LocalMux I__6196 (
            .O(N__32949),
            .I(N__32941));
    LocalMux I__6195 (
            .O(N__32946),
            .I(N__32941));
    Span4Mux_h I__6194 (
            .O(N__32941),
            .I(N__32936));
    InMux I__6193 (
            .O(N__32940),
            .I(N__32931));
    InMux I__6192 (
            .O(N__32939),
            .I(N__32931));
    Odrv4 I__6191 (
            .O(N__32936),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6190 (
            .O(N__32931),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__6189 (
            .O(N__32926),
            .I(N__32923));
    InMux I__6188 (
            .O(N__32923),
            .I(N__32920));
    LocalMux I__6187 (
            .O(N__32920),
            .I(N__32917));
    Span4Mux_v I__6186 (
            .O(N__32917),
            .I(N__32914));
    Span4Mux_v I__6185 (
            .O(N__32914),
            .I(N__32911));
    Span4Mux_v I__6184 (
            .O(N__32911),
            .I(N__32908));
    Odrv4 I__6183 (
            .O(N__32908),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__6182 (
            .O(N__32905),
            .I(N__32902));
    LocalMux I__6181 (
            .O(N__32902),
            .I(N__32899));
    Span4Mux_h I__6180 (
            .O(N__32899),
            .I(N__32894));
    InMux I__6179 (
            .O(N__32898),
            .I(N__32891));
    InMux I__6178 (
            .O(N__32897),
            .I(N__32888));
    Odrv4 I__6177 (
            .O(N__32894),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__6176 (
            .O(N__32891),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__6175 (
            .O(N__32888),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CEMux I__6174 (
            .O(N__32881),
            .I(N__32857));
    CEMux I__6173 (
            .O(N__32880),
            .I(N__32857));
    CEMux I__6172 (
            .O(N__32879),
            .I(N__32857));
    CEMux I__6171 (
            .O(N__32878),
            .I(N__32857));
    CEMux I__6170 (
            .O(N__32877),
            .I(N__32857));
    CEMux I__6169 (
            .O(N__32876),
            .I(N__32857));
    CEMux I__6168 (
            .O(N__32875),
            .I(N__32857));
    CEMux I__6167 (
            .O(N__32874),
            .I(N__32857));
    GlobalMux I__6166 (
            .O(N__32857),
            .I(N__32854));
    gio2CtrlBuf I__6165 (
            .O(N__32854),
            .I(\current_shift_inst.timer_s1.N_161_i_g ));
    InMux I__6164 (
            .O(N__32851),
            .I(N__32848));
    LocalMux I__6163 (
            .O(N__32848),
            .I(N__32845));
    Span4Mux_v I__6162 (
            .O(N__32845),
            .I(N__32842));
    Odrv4 I__6161 (
            .O(N__32842),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__6160 (
            .O(N__32839),
            .I(N__32835));
    InMux I__6159 (
            .O(N__32838),
            .I(N__32829));
    InMux I__6158 (
            .O(N__32835),
            .I(N__32829));
    InMux I__6157 (
            .O(N__32834),
            .I(N__32826));
    LocalMux I__6156 (
            .O(N__32829),
            .I(N__32823));
    LocalMux I__6155 (
            .O(N__32826),
            .I(N__32819));
    Span12Mux_h I__6154 (
            .O(N__32823),
            .I(N__32816));
    InMux I__6153 (
            .O(N__32822),
            .I(N__32813));
    Span4Mux_v I__6152 (
            .O(N__32819),
            .I(N__32810));
    Odrv12 I__6151 (
            .O(N__32816),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__6150 (
            .O(N__32813),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__6149 (
            .O(N__32810),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__6148 (
            .O(N__32803),
            .I(N__32800));
    InMux I__6147 (
            .O(N__32800),
            .I(N__32797));
    LocalMux I__6146 (
            .O(N__32797),
            .I(N__32794));
    Span4Mux_v I__6145 (
            .O(N__32794),
            .I(N__32791));
    Odrv4 I__6144 (
            .O(N__32791),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__6143 (
            .O(N__32788),
            .I(N__32772));
    InMux I__6142 (
            .O(N__32787),
            .I(N__32769));
    InMux I__6141 (
            .O(N__32786),
            .I(N__32764));
    InMux I__6140 (
            .O(N__32785),
            .I(N__32764));
    InMux I__6139 (
            .O(N__32784),
            .I(N__32748));
    InMux I__6138 (
            .O(N__32783),
            .I(N__32748));
    InMux I__6137 (
            .O(N__32782),
            .I(N__32748));
    InMux I__6136 (
            .O(N__32781),
            .I(N__32748));
    InMux I__6135 (
            .O(N__32780),
            .I(N__32748));
    InMux I__6134 (
            .O(N__32779),
            .I(N__32748));
    InMux I__6133 (
            .O(N__32778),
            .I(N__32745));
    InMux I__6132 (
            .O(N__32777),
            .I(N__32740));
    InMux I__6131 (
            .O(N__32776),
            .I(N__32735));
    InMux I__6130 (
            .O(N__32775),
            .I(N__32735));
    LocalMux I__6129 (
            .O(N__32772),
            .I(N__32728));
    LocalMux I__6128 (
            .O(N__32769),
            .I(N__32728));
    LocalMux I__6127 (
            .O(N__32764),
            .I(N__32728));
    InMux I__6126 (
            .O(N__32763),
            .I(N__32721));
    InMux I__6125 (
            .O(N__32762),
            .I(N__32721));
    InMux I__6124 (
            .O(N__32761),
            .I(N__32721));
    LocalMux I__6123 (
            .O(N__32748),
            .I(N__32718));
    LocalMux I__6122 (
            .O(N__32745),
            .I(N__32715));
    InMux I__6121 (
            .O(N__32744),
            .I(N__32710));
    InMux I__6120 (
            .O(N__32743),
            .I(N__32710));
    LocalMux I__6119 (
            .O(N__32740),
            .I(N__32705));
    LocalMux I__6118 (
            .O(N__32735),
            .I(N__32701));
    Span4Mux_v I__6117 (
            .O(N__32728),
            .I(N__32690));
    LocalMux I__6116 (
            .O(N__32721),
            .I(N__32690));
    Span4Mux_h I__6115 (
            .O(N__32718),
            .I(N__32690));
    Span4Mux_h I__6114 (
            .O(N__32715),
            .I(N__32690));
    LocalMux I__6113 (
            .O(N__32710),
            .I(N__32690));
    InMux I__6112 (
            .O(N__32709),
            .I(N__32685));
    InMux I__6111 (
            .O(N__32708),
            .I(N__32685));
    Span4Mux_h I__6110 (
            .O(N__32705),
            .I(N__32679));
    InMux I__6109 (
            .O(N__32704),
            .I(N__32676));
    Span4Mux_v I__6108 (
            .O(N__32701),
            .I(N__32673));
    Span4Mux_v I__6107 (
            .O(N__32690),
            .I(N__32668));
    LocalMux I__6106 (
            .O(N__32685),
            .I(N__32668));
    InMux I__6105 (
            .O(N__32684),
            .I(N__32665));
    InMux I__6104 (
            .O(N__32683),
            .I(N__32660));
    InMux I__6103 (
            .O(N__32682),
            .I(N__32660));
    Odrv4 I__6102 (
            .O(N__32679),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__6101 (
            .O(N__32676),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__6100 (
            .O(N__32673),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__6099 (
            .O(N__32668),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__6098 (
            .O(N__32665),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__6097 (
            .O(N__32660),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__6096 (
            .O(N__32647),
            .I(N__32644));
    InMux I__6095 (
            .O(N__32644),
            .I(N__32635));
    InMux I__6094 (
            .O(N__32643),
            .I(N__32635));
    InMux I__6093 (
            .O(N__32642),
            .I(N__32635));
    LocalMux I__6092 (
            .O(N__32635),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__6091 (
            .O(N__32632),
            .I(N__32620));
    InMux I__6090 (
            .O(N__32631),
            .I(N__32620));
    InMux I__6089 (
            .O(N__32630),
            .I(N__32620));
    InMux I__6088 (
            .O(N__32629),
            .I(N__32620));
    LocalMux I__6087 (
            .O(N__32620),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__6086 (
            .O(N__32617),
            .I(N__32614));
    InMux I__6085 (
            .O(N__32614),
            .I(N__32611));
    LocalMux I__6084 (
            .O(N__32611),
            .I(N__32608));
    Span4Mux_v I__6083 (
            .O(N__32608),
            .I(N__32605));
    Span4Mux_v I__6082 (
            .O(N__32605),
            .I(N__32602));
    Odrv4 I__6081 (
            .O(N__32602),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__6080 (
            .O(N__32599),
            .I(N__32593));
    CascadeMux I__6079 (
            .O(N__32598),
            .I(N__32590));
    InMux I__6078 (
            .O(N__32597),
            .I(N__32585));
    InMux I__6077 (
            .O(N__32596),
            .I(N__32585));
    InMux I__6076 (
            .O(N__32593),
            .I(N__32581));
    InMux I__6075 (
            .O(N__32590),
            .I(N__32578));
    LocalMux I__6074 (
            .O(N__32585),
            .I(N__32575));
    InMux I__6073 (
            .O(N__32584),
            .I(N__32572));
    LocalMux I__6072 (
            .O(N__32581),
            .I(N__32569));
    LocalMux I__6071 (
            .O(N__32578),
            .I(N__32566));
    Span4Mux_h I__6070 (
            .O(N__32575),
            .I(N__32563));
    LocalMux I__6069 (
            .O(N__32572),
            .I(N__32560));
    Span12Mux_s10_v I__6068 (
            .O(N__32569),
            .I(N__32557));
    Span4Mux_h I__6067 (
            .O(N__32566),
            .I(N__32552));
    Span4Mux_v I__6066 (
            .O(N__32563),
            .I(N__32552));
    Span4Mux_h I__6065 (
            .O(N__32560),
            .I(N__32549));
    Odrv12 I__6064 (
            .O(N__32557),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__6063 (
            .O(N__32552),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__6062 (
            .O(N__32549),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__6061 (
            .O(N__32542),
            .I(N__32538));
    InMux I__6060 (
            .O(N__32541),
            .I(N__32535));
    LocalMux I__6059 (
            .O(N__32538),
            .I(N__32529));
    LocalMux I__6058 (
            .O(N__32535),
            .I(N__32529));
    InMux I__6057 (
            .O(N__32534),
            .I(N__32526));
    Span4Mux_v I__6056 (
            .O(N__32529),
            .I(N__32523));
    LocalMux I__6055 (
            .O(N__32526),
            .I(N__32520));
    Span4Mux_v I__6054 (
            .O(N__32523),
            .I(N__32517));
    Odrv4 I__6053 (
            .O(N__32520),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__6052 (
            .O(N__32517),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__6051 (
            .O(N__32512),
            .I(N__32509));
    InMux I__6050 (
            .O(N__32509),
            .I(N__32506));
    LocalMux I__6049 (
            .O(N__32506),
            .I(N__32503));
    Span4Mux_h I__6048 (
            .O(N__32503),
            .I(N__32500));
    Odrv4 I__6047 (
            .O(N__32500),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__6046 (
            .O(N__32497),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__6045 (
            .O(N__32494),
            .I(N__32491));
    LocalMux I__6044 (
            .O(N__32491),
            .I(N__32485));
    InMux I__6043 (
            .O(N__32490),
            .I(N__32482));
    InMux I__6042 (
            .O(N__32489),
            .I(N__32477));
    InMux I__6041 (
            .O(N__32488),
            .I(N__32477));
    Odrv12 I__6040 (
            .O(N__32485),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__6039 (
            .O(N__32482),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__6038 (
            .O(N__32477),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    CascadeMux I__6037 (
            .O(N__32470),
            .I(N__32466));
    InMux I__6036 (
            .O(N__32469),
            .I(N__32463));
    InMux I__6035 (
            .O(N__32466),
            .I(N__32459));
    LocalMux I__6034 (
            .O(N__32463),
            .I(N__32456));
    InMux I__6033 (
            .O(N__32462),
            .I(N__32453));
    LocalMux I__6032 (
            .O(N__32459),
            .I(N__32450));
    Span4Mux_h I__6031 (
            .O(N__32456),
            .I(N__32447));
    LocalMux I__6030 (
            .O(N__32453),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__6029 (
            .O(N__32450),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__6028 (
            .O(N__32447),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__6027 (
            .O(N__32440),
            .I(N__32437));
    LocalMux I__6026 (
            .O(N__32437),
            .I(N__32434));
    Span4Mux_h I__6025 (
            .O(N__32434),
            .I(N__32431));
    Odrv4 I__6024 (
            .O(N__32431),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    CascadeMux I__6023 (
            .O(N__32428),
            .I(N__32425));
    InMux I__6022 (
            .O(N__32425),
            .I(N__32421));
    InMux I__6021 (
            .O(N__32424),
            .I(N__32418));
    LocalMux I__6020 (
            .O(N__32421),
            .I(N__32415));
    LocalMux I__6019 (
            .O(N__32418),
            .I(N__32412));
    Span4Mux_v I__6018 (
            .O(N__32415),
            .I(N__32408));
    Sp12to4 I__6017 (
            .O(N__32412),
            .I(N__32405));
    InMux I__6016 (
            .O(N__32411),
            .I(N__32402));
    Odrv4 I__6015 (
            .O(N__32408),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv12 I__6014 (
            .O(N__32405),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__6013 (
            .O(N__32402),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__6012 (
            .O(N__32395),
            .I(N__32392));
    InMux I__6011 (
            .O(N__32392),
            .I(N__32388));
    InMux I__6010 (
            .O(N__32391),
            .I(N__32385));
    LocalMux I__6009 (
            .O(N__32388),
            .I(N__32382));
    LocalMux I__6008 (
            .O(N__32385),
            .I(N__32377));
    Span4Mux_v I__6007 (
            .O(N__32382),
            .I(N__32377));
    Span4Mux_v I__6006 (
            .O(N__32377),
            .I(N__32373));
    InMux I__6005 (
            .O(N__32376),
            .I(N__32370));
    Span4Mux_h I__6004 (
            .O(N__32373),
            .I(N__32366));
    LocalMux I__6003 (
            .O(N__32370),
            .I(N__32363));
    InMux I__6002 (
            .O(N__32369),
            .I(N__32360));
    Odrv4 I__6001 (
            .O(N__32366),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__6000 (
            .O(N__32363),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__5999 (
            .O(N__32360),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__5998 (
            .O(N__32353),
            .I(N__32350));
    LocalMux I__5997 (
            .O(N__32350),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__5996 (
            .O(N__32347),
            .I(N__32344));
    LocalMux I__5995 (
            .O(N__32344),
            .I(N__32341));
    Span4Mux_h I__5994 (
            .O(N__32341),
            .I(N__32338));
    Span4Mux_v I__5993 (
            .O(N__32338),
            .I(N__32335));
    Odrv4 I__5992 (
            .O(N__32335),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__5991 (
            .O(N__32332),
            .I(N__32329));
    LocalMux I__5990 (
            .O(N__32329),
            .I(N__32326));
    Span4Mux_h I__5989 (
            .O(N__32326),
            .I(N__32323));
    Odrv4 I__5988 (
            .O(N__32323),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__5987 (
            .O(N__32320),
            .I(N__32317));
    LocalMux I__5986 (
            .O(N__32317),
            .I(N__32314));
    Span4Mux_h I__5985 (
            .O(N__32314),
            .I(N__32311));
    Span4Mux_v I__5984 (
            .O(N__32311),
            .I(N__32308));
    Odrv4 I__5983 (
            .O(N__32308),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__5982 (
            .O(N__32305),
            .I(N__32301));
    InMux I__5981 (
            .O(N__32304),
            .I(N__32295));
    InMux I__5980 (
            .O(N__32301),
            .I(N__32295));
    InMux I__5979 (
            .O(N__32300),
            .I(N__32292));
    LocalMux I__5978 (
            .O(N__32295),
            .I(N__32287));
    LocalMux I__5977 (
            .O(N__32292),
            .I(N__32287));
    Span4Mux_h I__5976 (
            .O(N__32287),
            .I(N__32283));
    InMux I__5975 (
            .O(N__32286),
            .I(N__32280));
    Odrv4 I__5974 (
            .O(N__32283),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__5973 (
            .O(N__32280),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__5972 (
            .O(N__32275),
            .I(N__32266));
    InMux I__5971 (
            .O(N__32274),
            .I(N__32266));
    InMux I__5970 (
            .O(N__32273),
            .I(N__32266));
    LocalMux I__5969 (
            .O(N__32266),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__5968 (
            .O(N__32263),
            .I(N__32260));
    LocalMux I__5967 (
            .O(N__32260),
            .I(N__32257));
    Span4Mux_h I__5966 (
            .O(N__32257),
            .I(N__32254));
    Span4Mux_v I__5965 (
            .O(N__32254),
            .I(N__32251));
    Odrv4 I__5964 (
            .O(N__32251),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__5963 (
            .O(N__32248),
            .I(N__32244));
    CascadeMux I__5962 (
            .O(N__32247),
            .I(N__32241));
    LocalMux I__5961 (
            .O(N__32244),
            .I(N__32238));
    InMux I__5960 (
            .O(N__32241),
            .I(N__32234));
    Span4Mux_h I__5959 (
            .O(N__32238),
            .I(N__32231));
    InMux I__5958 (
            .O(N__32237),
            .I(N__32228));
    LocalMux I__5957 (
            .O(N__32234),
            .I(N__32225));
    Odrv4 I__5956 (
            .O(N__32231),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__5955 (
            .O(N__32228),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__5954 (
            .O(N__32225),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__5953 (
            .O(N__32218),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__5952 (
            .O(N__32215),
            .I(N__32212));
    InMux I__5951 (
            .O(N__32212),
            .I(N__32208));
    InMux I__5950 (
            .O(N__32211),
            .I(N__32205));
    LocalMux I__5949 (
            .O(N__32208),
            .I(N__32202));
    LocalMux I__5948 (
            .O(N__32205),
            .I(N__32199));
    Span4Mux_h I__5947 (
            .O(N__32202),
            .I(N__32196));
    Span4Mux_h I__5946 (
            .O(N__32199),
            .I(N__32191));
    Span4Mux_v I__5945 (
            .O(N__32196),
            .I(N__32191));
    Odrv4 I__5944 (
            .O(N__32191),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__5943 (
            .O(N__32188),
            .I(N__32185));
    LocalMux I__5942 (
            .O(N__32185),
            .I(N__32180));
    InMux I__5941 (
            .O(N__32184),
            .I(N__32177));
    InMux I__5940 (
            .O(N__32183),
            .I(N__32174));
    Span4Mux_h I__5939 (
            .O(N__32180),
            .I(N__32171));
    LocalMux I__5938 (
            .O(N__32177),
            .I(N__32168));
    LocalMux I__5937 (
            .O(N__32174),
            .I(N__32165));
    Span4Mux_v I__5936 (
            .O(N__32171),
            .I(N__32160));
    Span4Mux_h I__5935 (
            .O(N__32168),
            .I(N__32160));
    Odrv4 I__5934 (
            .O(N__32165),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__5933 (
            .O(N__32160),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CascadeMux I__5932 (
            .O(N__32155),
            .I(N__32152));
    InMux I__5931 (
            .O(N__32152),
            .I(N__32148));
    CascadeMux I__5930 (
            .O(N__32151),
            .I(N__32145));
    LocalMux I__5929 (
            .O(N__32148),
            .I(N__32142));
    InMux I__5928 (
            .O(N__32145),
            .I(N__32139));
    Span4Mux_h I__5927 (
            .O(N__32142),
            .I(N__32133));
    LocalMux I__5926 (
            .O(N__32139),
            .I(N__32133));
    InMux I__5925 (
            .O(N__32138),
            .I(N__32130));
    Span4Mux_v I__5924 (
            .O(N__32133),
            .I(N__32126));
    LocalMux I__5923 (
            .O(N__32130),
            .I(N__32123));
    InMux I__5922 (
            .O(N__32129),
            .I(N__32120));
    Odrv4 I__5921 (
            .O(N__32126),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__5920 (
            .O(N__32123),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__5919 (
            .O(N__32120),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__5918 (
            .O(N__32113),
            .I(N__32108));
    InMux I__5917 (
            .O(N__32112),
            .I(N__32105));
    InMux I__5916 (
            .O(N__32111),
            .I(N__32102));
    LocalMux I__5915 (
            .O(N__32108),
            .I(N__32099));
    LocalMux I__5914 (
            .O(N__32105),
            .I(N__32096));
    LocalMux I__5913 (
            .O(N__32102),
            .I(N__32093));
    Span4Mux_v I__5912 (
            .O(N__32099),
            .I(N__32090));
    Odrv12 I__5911 (
            .O(N__32096),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__5910 (
            .O(N__32093),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__5909 (
            .O(N__32090),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__5908 (
            .O(N__32083),
            .I(N__32080));
    InMux I__5907 (
            .O(N__32080),
            .I(N__32077));
    LocalMux I__5906 (
            .O(N__32077),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    CascadeMux I__5905 (
            .O(N__32074),
            .I(N__32071));
    InMux I__5904 (
            .O(N__32071),
            .I(N__32068));
    LocalMux I__5903 (
            .O(N__32068),
            .I(N__32064));
    InMux I__5902 (
            .O(N__32067),
            .I(N__32061));
    Span4Mux_v I__5901 (
            .O(N__32064),
            .I(N__32056));
    LocalMux I__5900 (
            .O(N__32061),
            .I(N__32056));
    Span4Mux_v I__5899 (
            .O(N__32056),
            .I(N__32053));
    Span4Mux_h I__5898 (
            .O(N__32053),
            .I(N__32049));
    InMux I__5897 (
            .O(N__32052),
            .I(N__32046));
    Odrv4 I__5896 (
            .O(N__32049),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__5895 (
            .O(N__32046),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__5894 (
            .O(N__32041),
            .I(N__32038));
    InMux I__5893 (
            .O(N__32038),
            .I(N__32034));
    InMux I__5892 (
            .O(N__32037),
            .I(N__32031));
    LocalMux I__5891 (
            .O(N__32034),
            .I(N__32027));
    LocalMux I__5890 (
            .O(N__32031),
            .I(N__32024));
    InMux I__5889 (
            .O(N__32030),
            .I(N__32020));
    Span4Mux_h I__5888 (
            .O(N__32027),
            .I(N__32017));
    Span12Mux_v I__5887 (
            .O(N__32024),
            .I(N__32014));
    InMux I__5886 (
            .O(N__32023),
            .I(N__32011));
    LocalMux I__5885 (
            .O(N__32020),
            .I(N__32008));
    Odrv4 I__5884 (
            .O(N__32017),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__5883 (
            .O(N__32014),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__5882 (
            .O(N__32011),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__5881 (
            .O(N__32008),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    CascadeMux I__5880 (
            .O(N__31999),
            .I(N__31996));
    InMux I__5879 (
            .O(N__31996),
            .I(N__31993));
    LocalMux I__5878 (
            .O(N__31993),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__5877 (
            .O(N__31990),
            .I(N__31986));
    InMux I__5876 (
            .O(N__31989),
            .I(N__31982));
    InMux I__5875 (
            .O(N__31986),
            .I(N__31979));
    InMux I__5874 (
            .O(N__31985),
            .I(N__31976));
    LocalMux I__5873 (
            .O(N__31982),
            .I(N__31973));
    LocalMux I__5872 (
            .O(N__31979),
            .I(N__31970));
    LocalMux I__5871 (
            .O(N__31976),
            .I(N__31965));
    Span4Mux_h I__5870 (
            .O(N__31973),
            .I(N__31965));
    Odrv4 I__5869 (
            .O(N__31970),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__5868 (
            .O(N__31965),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__5867 (
            .O(N__31960),
            .I(N__31957));
    LocalMux I__5866 (
            .O(N__31957),
            .I(N__31953));
    CascadeMux I__5865 (
            .O(N__31956),
            .I(N__31949));
    Span4Mux_v I__5864 (
            .O(N__31953),
            .I(N__31946));
    InMux I__5863 (
            .O(N__31952),
            .I(N__31943));
    InMux I__5862 (
            .O(N__31949),
            .I(N__31939));
    Span4Mux_h I__5861 (
            .O(N__31946),
            .I(N__31934));
    LocalMux I__5860 (
            .O(N__31943),
            .I(N__31934));
    InMux I__5859 (
            .O(N__31942),
            .I(N__31931));
    LocalMux I__5858 (
            .O(N__31939),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__5857 (
            .O(N__31934),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__5856 (
            .O(N__31931),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    CascadeMux I__5855 (
            .O(N__31924),
            .I(N__31921));
    InMux I__5854 (
            .O(N__31921),
            .I(N__31918));
    LocalMux I__5853 (
            .O(N__31918),
            .I(N__31915));
    Span4Mux_h I__5852 (
            .O(N__31915),
            .I(N__31912));
    Span4Mux_h I__5851 (
            .O(N__31912),
            .I(N__31909));
    Odrv4 I__5850 (
            .O(N__31909),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    CascadeMux I__5849 (
            .O(N__31906),
            .I(N__31903));
    InMux I__5848 (
            .O(N__31903),
            .I(N__31900));
    LocalMux I__5847 (
            .O(N__31900),
            .I(N__31897));
    Odrv4 I__5846 (
            .O(N__31897),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__5845 (
            .O(N__31894),
            .I(N__31891));
    LocalMux I__5844 (
            .O(N__31891),
            .I(N__31888));
    Span4Mux_v I__5843 (
            .O(N__31888),
            .I(N__31883));
    InMux I__5842 (
            .O(N__31887),
            .I(N__31878));
    InMux I__5841 (
            .O(N__31886),
            .I(N__31878));
    Odrv4 I__5840 (
            .O(N__31883),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__5839 (
            .O(N__31878),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__5838 (
            .O(N__31873),
            .I(N__31869));
    CascadeMux I__5837 (
            .O(N__31872),
            .I(N__31866));
    InMux I__5836 (
            .O(N__31869),
            .I(N__31862));
    InMux I__5835 (
            .O(N__31866),
            .I(N__31857));
    InMux I__5834 (
            .O(N__31865),
            .I(N__31857));
    LocalMux I__5833 (
            .O(N__31862),
            .I(N__31854));
    LocalMux I__5832 (
            .O(N__31857),
            .I(N__31851));
    Span12Mux_v I__5831 (
            .O(N__31854),
            .I(N__31847));
    Span4Mux_h I__5830 (
            .O(N__31851),
            .I(N__31844));
    InMux I__5829 (
            .O(N__31850),
            .I(N__31841));
    Odrv12 I__5828 (
            .O(N__31847),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__5827 (
            .O(N__31844),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__5826 (
            .O(N__31841),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    CascadeMux I__5825 (
            .O(N__31834),
            .I(N__31831));
    InMux I__5824 (
            .O(N__31831),
            .I(N__31828));
    LocalMux I__5823 (
            .O(N__31828),
            .I(N__31825));
    Span4Mux_h I__5822 (
            .O(N__31825),
            .I(N__31822));
    Odrv4 I__5821 (
            .O(N__31822),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__5820 (
            .O(N__31819),
            .I(N__31815));
    InMux I__5819 (
            .O(N__31818),
            .I(N__31811));
    LocalMux I__5818 (
            .O(N__31815),
            .I(N__31808));
    CascadeMux I__5817 (
            .O(N__31814),
            .I(N__31805));
    LocalMux I__5816 (
            .O(N__31811),
            .I(N__31802));
    Span4Mux_v I__5815 (
            .O(N__31808),
            .I(N__31799));
    InMux I__5814 (
            .O(N__31805),
            .I(N__31796));
    Span4Mux_v I__5813 (
            .O(N__31802),
            .I(N__31793));
    Odrv4 I__5812 (
            .O(N__31799),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__5811 (
            .O(N__31796),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__5810 (
            .O(N__31793),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__5809 (
            .O(N__31786),
            .I(N__31783));
    LocalMux I__5808 (
            .O(N__31783),
            .I(N__31779));
    CascadeMux I__5807 (
            .O(N__31782),
            .I(N__31775));
    Span4Mux_v I__5806 (
            .O(N__31779),
            .I(N__31772));
    InMux I__5805 (
            .O(N__31778),
            .I(N__31769));
    InMux I__5804 (
            .O(N__31775),
            .I(N__31766));
    Span4Mux_v I__5803 (
            .O(N__31772),
            .I(N__31761));
    LocalMux I__5802 (
            .O(N__31769),
            .I(N__31761));
    LocalMux I__5801 (
            .O(N__31766),
            .I(N__31757));
    Span4Mux_h I__5800 (
            .O(N__31761),
            .I(N__31754));
    InMux I__5799 (
            .O(N__31760),
            .I(N__31751));
    Odrv12 I__5798 (
            .O(N__31757),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__5797 (
            .O(N__31754),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__5796 (
            .O(N__31751),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__5795 (
            .O(N__31744),
            .I(N__31741));
    LocalMux I__5794 (
            .O(N__31741),
            .I(N__31738));
    Span4Mux_h I__5793 (
            .O(N__31738),
            .I(N__31735));
    Span4Mux_v I__5792 (
            .O(N__31735),
            .I(N__31732));
    Odrv4 I__5791 (
            .O(N__31732),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    CascadeMux I__5790 (
            .O(N__31729),
            .I(N__31726));
    InMux I__5789 (
            .O(N__31726),
            .I(N__31723));
    LocalMux I__5788 (
            .O(N__31723),
            .I(N__31719));
    CascadeMux I__5787 (
            .O(N__31722),
            .I(N__31716));
    Span4Mux_h I__5786 (
            .O(N__31719),
            .I(N__31712));
    InMux I__5785 (
            .O(N__31716),
            .I(N__31709));
    InMux I__5784 (
            .O(N__31715),
            .I(N__31706));
    Span4Mux_v I__5783 (
            .O(N__31712),
            .I(N__31702));
    LocalMux I__5782 (
            .O(N__31709),
            .I(N__31699));
    LocalMux I__5781 (
            .O(N__31706),
            .I(N__31696));
    InMux I__5780 (
            .O(N__31705),
            .I(N__31693));
    Odrv4 I__5779 (
            .O(N__31702),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv12 I__5778 (
            .O(N__31699),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__5777 (
            .O(N__31696),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__5776 (
            .O(N__31693),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__5775 (
            .O(N__31684),
            .I(N__31679));
    InMux I__5774 (
            .O(N__31683),
            .I(N__31676));
    InMux I__5773 (
            .O(N__31682),
            .I(N__31673));
    LocalMux I__5772 (
            .O(N__31679),
            .I(N__31670));
    LocalMux I__5771 (
            .O(N__31676),
            .I(N__31667));
    LocalMux I__5770 (
            .O(N__31673),
            .I(N__31664));
    Span4Mux_v I__5769 (
            .O(N__31670),
            .I(N__31661));
    Odrv12 I__5768 (
            .O(N__31667),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__5767 (
            .O(N__31664),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__5766 (
            .O(N__31661),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__5765 (
            .O(N__31654),
            .I(N__31651));
    InMux I__5764 (
            .O(N__31651),
            .I(N__31648));
    LocalMux I__5763 (
            .O(N__31648),
            .I(N__31645));
    Odrv4 I__5762 (
            .O(N__31645),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    CascadeMux I__5761 (
            .O(N__31642),
            .I(N__31638));
    InMux I__5760 (
            .O(N__31641),
            .I(N__31635));
    InMux I__5759 (
            .O(N__31638),
            .I(N__31632));
    LocalMux I__5758 (
            .O(N__31635),
            .I(N__31629));
    LocalMux I__5757 (
            .O(N__31632),
            .I(N__31623));
    Span4Mux_v I__5756 (
            .O(N__31629),
            .I(N__31623));
    InMux I__5755 (
            .O(N__31628),
            .I(N__31620));
    Span4Mux_v I__5754 (
            .O(N__31623),
            .I(N__31616));
    LocalMux I__5753 (
            .O(N__31620),
            .I(N__31613));
    InMux I__5752 (
            .O(N__31619),
            .I(N__31610));
    Odrv4 I__5751 (
            .O(N__31616),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__5750 (
            .O(N__31613),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__5749 (
            .O(N__31610),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    CascadeMux I__5748 (
            .O(N__31603),
            .I(N__31600));
    InMux I__5747 (
            .O(N__31600),
            .I(N__31595));
    InMux I__5746 (
            .O(N__31599),
            .I(N__31592));
    InMux I__5745 (
            .O(N__31598),
            .I(N__31589));
    LocalMux I__5744 (
            .O(N__31595),
            .I(N__31586));
    LocalMux I__5743 (
            .O(N__31592),
            .I(N__31583));
    LocalMux I__5742 (
            .O(N__31589),
            .I(N__31580));
    Span4Mux_v I__5741 (
            .O(N__31586),
            .I(N__31575));
    Span4Mux_v I__5740 (
            .O(N__31583),
            .I(N__31575));
    Odrv4 I__5739 (
            .O(N__31580),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__5738 (
            .O(N__31575),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__5737 (
            .O(N__31570),
            .I(N__31567));
    LocalMux I__5736 (
            .O(N__31567),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    CascadeMux I__5735 (
            .O(N__31564),
            .I(N__31561));
    InMux I__5734 (
            .O(N__31561),
            .I(N__31558));
    LocalMux I__5733 (
            .O(N__31558),
            .I(N__31554));
    InMux I__5732 (
            .O(N__31557),
            .I(N__31551));
    Span4Mux_v I__5731 (
            .O(N__31554),
            .I(N__31547));
    LocalMux I__5730 (
            .O(N__31551),
            .I(N__31544));
    InMux I__5729 (
            .O(N__31550),
            .I(N__31541));
    Span4Mux_h I__5728 (
            .O(N__31547),
            .I(N__31538));
    Span4Mux_v I__5727 (
            .O(N__31544),
            .I(N__31535));
    LocalMux I__5726 (
            .O(N__31541),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__5725 (
            .O(N__31538),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__5724 (
            .O(N__31535),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__5723 (
            .O(N__31528),
            .I(N__31524));
    CascadeMux I__5722 (
            .O(N__31527),
            .I(N__31520));
    LocalMux I__5721 (
            .O(N__31524),
            .I(N__31516));
    InMux I__5720 (
            .O(N__31523),
            .I(N__31513));
    InMux I__5719 (
            .O(N__31520),
            .I(N__31508));
    InMux I__5718 (
            .O(N__31519),
            .I(N__31508));
    Span4Mux_h I__5717 (
            .O(N__31516),
            .I(N__31503));
    LocalMux I__5716 (
            .O(N__31513),
            .I(N__31503));
    LocalMux I__5715 (
            .O(N__31508),
            .I(N__31500));
    Odrv4 I__5714 (
            .O(N__31503),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__5713 (
            .O(N__31500),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    CascadeMux I__5712 (
            .O(N__31495),
            .I(N__31492));
    InMux I__5711 (
            .O(N__31492),
            .I(N__31489));
    LocalMux I__5710 (
            .O(N__31489),
            .I(N__31486));
    Odrv4 I__5709 (
            .O(N__31486),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__5708 (
            .O(N__31483),
            .I(N__31479));
    CascadeMux I__5707 (
            .O(N__31482),
            .I(N__31476));
    InMux I__5706 (
            .O(N__31479),
            .I(N__31472));
    InMux I__5705 (
            .O(N__31476),
            .I(N__31469));
    InMux I__5704 (
            .O(N__31475),
            .I(N__31466));
    LocalMux I__5703 (
            .O(N__31472),
            .I(N__31461));
    LocalMux I__5702 (
            .O(N__31469),
            .I(N__31461));
    LocalMux I__5701 (
            .O(N__31466),
            .I(N__31458));
    Span4Mux_v I__5700 (
            .O(N__31461),
            .I(N__31454));
    Span4Mux_v I__5699 (
            .O(N__31458),
            .I(N__31451));
    InMux I__5698 (
            .O(N__31457),
            .I(N__31448));
    Odrv4 I__5697 (
            .O(N__31454),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__5696 (
            .O(N__31451),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__5695 (
            .O(N__31448),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__5694 (
            .O(N__31441),
            .I(N__31438));
    LocalMux I__5693 (
            .O(N__31438),
            .I(N__31434));
    InMux I__5692 (
            .O(N__31437),
            .I(N__31431));
    Span4Mux_h I__5691 (
            .O(N__31434),
            .I(N__31425));
    LocalMux I__5690 (
            .O(N__31431),
            .I(N__31425));
    InMux I__5689 (
            .O(N__31430),
            .I(N__31422));
    Odrv4 I__5688 (
            .O(N__31425),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__5687 (
            .O(N__31422),
            .I(\current_shift_inst.un4_control_input1_3 ));
    CascadeMux I__5686 (
            .O(N__31417),
            .I(N__31414));
    InMux I__5685 (
            .O(N__31414),
            .I(N__31411));
    LocalMux I__5684 (
            .O(N__31411),
            .I(N__31408));
    Odrv4 I__5683 (
            .O(N__31408),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__5682 (
            .O(N__31405),
            .I(N__31402));
    InMux I__5681 (
            .O(N__31402),
            .I(N__31397));
    InMux I__5680 (
            .O(N__31401),
            .I(N__31394));
    InMux I__5679 (
            .O(N__31400),
            .I(N__31391));
    LocalMux I__5678 (
            .O(N__31397),
            .I(N__31388));
    LocalMux I__5677 (
            .O(N__31394),
            .I(N__31385));
    LocalMux I__5676 (
            .O(N__31391),
            .I(N__31382));
    Span4Mux_v I__5675 (
            .O(N__31388),
            .I(N__31379));
    Span4Mux_v I__5674 (
            .O(N__31385),
            .I(N__31376));
    Odrv12 I__5673 (
            .O(N__31382),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__5672 (
            .O(N__31379),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__5671 (
            .O(N__31376),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__5670 (
            .O(N__31369),
            .I(N__31366));
    InMux I__5669 (
            .O(N__31366),
            .I(N__31362));
    InMux I__5668 (
            .O(N__31365),
            .I(N__31359));
    LocalMux I__5667 (
            .O(N__31362),
            .I(N__31355));
    LocalMux I__5666 (
            .O(N__31359),
            .I(N__31352));
    InMux I__5665 (
            .O(N__31358),
            .I(N__31349));
    Span4Mux_h I__5664 (
            .O(N__31355),
            .I(N__31345));
    Span4Mux_v I__5663 (
            .O(N__31352),
            .I(N__31340));
    LocalMux I__5662 (
            .O(N__31349),
            .I(N__31340));
    InMux I__5661 (
            .O(N__31348),
            .I(N__31337));
    Span4Mux_v I__5660 (
            .O(N__31345),
            .I(N__31334));
    Span4Mux_h I__5659 (
            .O(N__31340),
            .I(N__31331));
    LocalMux I__5658 (
            .O(N__31337),
            .I(N__31328));
    Odrv4 I__5657 (
            .O(N__31334),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__5656 (
            .O(N__31331),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__5655 (
            .O(N__31328),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__5654 (
            .O(N__31321),
            .I(N__31318));
    LocalMux I__5653 (
            .O(N__31318),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__5652 (
            .O(N__31315),
            .I(N__31312));
    LocalMux I__5651 (
            .O(N__31312),
            .I(N__31309));
    Odrv4 I__5650 (
            .O(N__31309),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    InMux I__5649 (
            .O(N__31306),
            .I(N__31303));
    LocalMux I__5648 (
            .O(N__31303),
            .I(N__31298));
    InMux I__5647 (
            .O(N__31302),
            .I(N__31295));
    InMux I__5646 (
            .O(N__31301),
            .I(N__31292));
    Span4Mux_v I__5645 (
            .O(N__31298),
            .I(N__31287));
    LocalMux I__5644 (
            .O(N__31295),
            .I(N__31287));
    LocalMux I__5643 (
            .O(N__31292),
            .I(N__31283));
    Span4Mux_h I__5642 (
            .O(N__31287),
            .I(N__31280));
    InMux I__5641 (
            .O(N__31286),
            .I(N__31277));
    Odrv4 I__5640 (
            .O(N__31283),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__5639 (
            .O(N__31280),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__5638 (
            .O(N__31277),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__5637 (
            .O(N__31270),
            .I(N__31265));
    InMux I__5636 (
            .O(N__31269),
            .I(N__31262));
    CascadeMux I__5635 (
            .O(N__31268),
            .I(N__31259));
    LocalMux I__5634 (
            .O(N__31265),
            .I(N__31256));
    LocalMux I__5633 (
            .O(N__31262),
            .I(N__31253));
    InMux I__5632 (
            .O(N__31259),
            .I(N__31250));
    Span4Mux_v I__5631 (
            .O(N__31256),
            .I(N__31247));
    Span4Mux_v I__5630 (
            .O(N__31253),
            .I(N__31244));
    LocalMux I__5629 (
            .O(N__31250),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__5628 (
            .O(N__31247),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__5627 (
            .O(N__31244),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__5626 (
            .O(N__31237),
            .I(N__31234));
    InMux I__5625 (
            .O(N__31234),
            .I(N__31231));
    LocalMux I__5624 (
            .O(N__31231),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__5623 (
            .O(N__31228),
            .I(N__31223));
    InMux I__5622 (
            .O(N__31227),
            .I(N__31217));
    InMux I__5621 (
            .O(N__31226),
            .I(N__31217));
    LocalMux I__5620 (
            .O(N__31223),
            .I(N__31214));
    InMux I__5619 (
            .O(N__31222),
            .I(N__31211));
    LocalMux I__5618 (
            .O(N__31217),
            .I(N__31208));
    Odrv4 I__5617 (
            .O(N__31214),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__5616 (
            .O(N__31211),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__5615 (
            .O(N__31208),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__5614 (
            .O(N__31201),
            .I(N__31196));
    InMux I__5613 (
            .O(N__31200),
            .I(N__31193));
    CascadeMux I__5612 (
            .O(N__31199),
            .I(N__31190));
    LocalMux I__5611 (
            .O(N__31196),
            .I(N__31187));
    LocalMux I__5610 (
            .O(N__31193),
            .I(N__31184));
    InMux I__5609 (
            .O(N__31190),
            .I(N__31181));
    Odrv4 I__5608 (
            .O(N__31187),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__5607 (
            .O(N__31184),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__5606 (
            .O(N__31181),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__5605 (
            .O(N__31174),
            .I(N__31171));
    InMux I__5604 (
            .O(N__31171),
            .I(N__31168));
    LocalMux I__5603 (
            .O(N__31168),
            .I(N__31165));
    Odrv4 I__5602 (
            .O(N__31165),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__5601 (
            .O(N__31162),
            .I(N__31158));
    CascadeMux I__5600 (
            .O(N__31161),
            .I(N__31155));
    LocalMux I__5599 (
            .O(N__31158),
            .I(N__31152));
    InMux I__5598 (
            .O(N__31155),
            .I(N__31149));
    Span4Mux_h I__5597 (
            .O(N__31152),
            .I(N__31146));
    LocalMux I__5596 (
            .O(N__31149),
            .I(N__31143));
    Span4Mux_v I__5595 (
            .O(N__31146),
            .I(N__31138));
    Span4Mux_h I__5594 (
            .O(N__31143),
            .I(N__31135));
    InMux I__5593 (
            .O(N__31142),
            .I(N__31132));
    InMux I__5592 (
            .O(N__31141),
            .I(N__31129));
    Odrv4 I__5591 (
            .O(N__31138),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__5590 (
            .O(N__31135),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__5589 (
            .O(N__31132),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__5588 (
            .O(N__31129),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__5587 (
            .O(N__31120),
            .I(N__31116));
    InMux I__5586 (
            .O(N__31119),
            .I(N__31113));
    LocalMux I__5585 (
            .O(N__31116),
            .I(N__31110));
    LocalMux I__5584 (
            .O(N__31113),
            .I(N__31107));
    Span4Mux_h I__5583 (
            .O(N__31110),
            .I(N__31104));
    Span4Mux_h I__5582 (
            .O(N__31107),
            .I(N__31098));
    Span4Mux_v I__5581 (
            .O(N__31104),
            .I(N__31098));
    InMux I__5580 (
            .O(N__31103),
            .I(N__31095));
    Odrv4 I__5579 (
            .O(N__31098),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__5578 (
            .O(N__31095),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__5577 (
            .O(N__31090),
            .I(N__31087));
    LocalMux I__5576 (
            .O(N__31087),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__5575 (
            .O(N__31084),
            .I(N__31081));
    LocalMux I__5574 (
            .O(N__31081),
            .I(N__31076));
    InMux I__5573 (
            .O(N__31080),
            .I(N__31073));
    InMux I__5572 (
            .O(N__31079),
            .I(N__31069));
    Span4Mux_h I__5571 (
            .O(N__31076),
            .I(N__31064));
    LocalMux I__5570 (
            .O(N__31073),
            .I(N__31064));
    InMux I__5569 (
            .O(N__31072),
            .I(N__31061));
    LocalMux I__5568 (
            .O(N__31069),
            .I(N__31058));
    Span4Mux_v I__5567 (
            .O(N__31064),
            .I(N__31053));
    LocalMux I__5566 (
            .O(N__31061),
            .I(N__31053));
    Span4Mux_v I__5565 (
            .O(N__31058),
            .I(N__31050));
    Span4Mux_h I__5564 (
            .O(N__31053),
            .I(N__31047));
    Odrv4 I__5563 (
            .O(N__31050),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__5562 (
            .O(N__31047),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__5561 (
            .O(N__31042),
            .I(N__31039));
    LocalMux I__5560 (
            .O(N__31039),
            .I(N__31036));
    Sp12to4 I__5559 (
            .O(N__31036),
            .I(N__31033));
    Odrv12 I__5558 (
            .O(N__31033),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__5557 (
            .O(N__31030),
            .I(N__31026));
    InMux I__5556 (
            .O(N__31029),
            .I(N__31023));
    LocalMux I__5555 (
            .O(N__31026),
            .I(N__31020));
    LocalMux I__5554 (
            .O(N__31023),
            .I(N__31017));
    Span4Mux_h I__5553 (
            .O(N__31020),
            .I(N__31014));
    Span4Mux_s3_h I__5552 (
            .O(N__31017),
            .I(N__31011));
    Span4Mux_h I__5551 (
            .O(N__31014),
            .I(N__31008));
    Span4Mux_h I__5550 (
            .O(N__31011),
            .I(N__31005));
    Odrv4 I__5549 (
            .O(N__31008),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__5548 (
            .O(N__31005),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__5547 (
            .O(N__31000),
            .I(N__30997));
    LocalMux I__5546 (
            .O(N__30997),
            .I(N__30994));
    Span4Mux_h I__5545 (
            .O(N__30994),
            .I(N__30991));
    Odrv4 I__5544 (
            .O(N__30991),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    CascadeMux I__5543 (
            .O(N__30988),
            .I(N__30984));
    CascadeMux I__5542 (
            .O(N__30987),
            .I(N__30981));
    InMux I__5541 (
            .O(N__30984),
            .I(N__30976));
    InMux I__5540 (
            .O(N__30981),
            .I(N__30976));
    LocalMux I__5539 (
            .O(N__30976),
            .I(N__30973));
    Span4Mux_h I__5538 (
            .O(N__30973),
            .I(N__30968));
    InMux I__5537 (
            .O(N__30972),
            .I(N__30963));
    InMux I__5536 (
            .O(N__30971),
            .I(N__30963));
    Odrv4 I__5535 (
            .O(N__30968),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__5534 (
            .O(N__30963),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__5533 (
            .O(N__30958),
            .I(N__30952));
    InMux I__5532 (
            .O(N__30957),
            .I(N__30952));
    LocalMux I__5531 (
            .O(N__30952),
            .I(N__30949));
    Span4Mux_h I__5530 (
            .O(N__30949),
            .I(N__30945));
    InMux I__5529 (
            .O(N__30948),
            .I(N__30942));
    Odrv4 I__5528 (
            .O(N__30945),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__5527 (
            .O(N__30942),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__5526 (
            .O(N__30937),
            .I(N__30934));
    LocalMux I__5525 (
            .O(N__30934),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    CascadeMux I__5524 (
            .O(N__30931),
            .I(N__30928));
    InMux I__5523 (
            .O(N__30928),
            .I(N__30925));
    LocalMux I__5522 (
            .O(N__30925),
            .I(N__30922));
    Span4Mux_h I__5521 (
            .O(N__30922),
            .I(N__30919));
    Span4Mux_v I__5520 (
            .O(N__30919),
            .I(N__30916));
    Odrv4 I__5519 (
            .O(N__30916),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__5518 (
            .O(N__30913),
            .I(N__30909));
    InMux I__5517 (
            .O(N__30912),
            .I(N__30905));
    InMux I__5516 (
            .O(N__30909),
            .I(N__30902));
    InMux I__5515 (
            .O(N__30908),
            .I(N__30899));
    LocalMux I__5514 (
            .O(N__30905),
            .I(N__30896));
    LocalMux I__5513 (
            .O(N__30902),
            .I(N__30893));
    LocalMux I__5512 (
            .O(N__30899),
            .I(N__30890));
    Span4Mux_v I__5511 (
            .O(N__30896),
            .I(N__30885));
    Span4Mux_h I__5510 (
            .O(N__30893),
            .I(N__30885));
    Span4Mux_v I__5509 (
            .O(N__30890),
            .I(N__30882));
    Odrv4 I__5508 (
            .O(N__30885),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__5507 (
            .O(N__30882),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__5506 (
            .O(N__30877),
            .I(N__30874));
    InMux I__5505 (
            .O(N__30874),
            .I(N__30871));
    LocalMux I__5504 (
            .O(N__30871),
            .I(N__30868));
    Odrv4 I__5503 (
            .O(N__30868),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    CascadeMux I__5502 (
            .O(N__30865),
            .I(N__30861));
    CascadeMux I__5501 (
            .O(N__30864),
            .I(N__30858));
    InMux I__5500 (
            .O(N__30861),
            .I(N__30855));
    InMux I__5499 (
            .O(N__30858),
            .I(N__30851));
    LocalMux I__5498 (
            .O(N__30855),
            .I(N__30848));
    InMux I__5497 (
            .O(N__30854),
            .I(N__30845));
    LocalMux I__5496 (
            .O(N__30851),
            .I(N__30841));
    Span4Mux_h I__5495 (
            .O(N__30848),
            .I(N__30838));
    LocalMux I__5494 (
            .O(N__30845),
            .I(N__30835));
    InMux I__5493 (
            .O(N__30844),
            .I(N__30832));
    Span4Mux_h I__5492 (
            .O(N__30841),
            .I(N__30829));
    Span4Mux_v I__5491 (
            .O(N__30838),
            .I(N__30826));
    Span4Mux_v I__5490 (
            .O(N__30835),
            .I(N__30821));
    LocalMux I__5489 (
            .O(N__30832),
            .I(N__30821));
    Odrv4 I__5488 (
            .O(N__30829),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__5487 (
            .O(N__30826),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__5486 (
            .O(N__30821),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__5485 (
            .O(N__30814),
            .I(N__30810));
    InMux I__5484 (
            .O(N__30813),
            .I(N__30806));
    LocalMux I__5483 (
            .O(N__30810),
            .I(N__30803));
    InMux I__5482 (
            .O(N__30809),
            .I(N__30800));
    LocalMux I__5481 (
            .O(N__30806),
            .I(N__30797));
    Span4Mux_v I__5480 (
            .O(N__30803),
            .I(N__30792));
    LocalMux I__5479 (
            .O(N__30800),
            .I(N__30792));
    Span4Mux_v I__5478 (
            .O(N__30797),
            .I(N__30789));
    Span4Mux_v I__5477 (
            .O(N__30792),
            .I(N__30786));
    Odrv4 I__5476 (
            .O(N__30789),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__5475 (
            .O(N__30786),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__5474 (
            .O(N__30781),
            .I(N__30778));
    InMux I__5473 (
            .O(N__30778),
            .I(N__30775));
    LocalMux I__5472 (
            .O(N__30775),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    CascadeMux I__5471 (
            .O(N__30772),
            .I(N__30769));
    InMux I__5470 (
            .O(N__30769),
            .I(N__30765));
    CascadeMux I__5469 (
            .O(N__30768),
            .I(N__30762));
    LocalMux I__5468 (
            .O(N__30765),
            .I(N__30758));
    InMux I__5467 (
            .O(N__30762),
            .I(N__30755));
    InMux I__5466 (
            .O(N__30761),
            .I(N__30752));
    Span4Mux_h I__5465 (
            .O(N__30758),
            .I(N__30748));
    LocalMux I__5464 (
            .O(N__30755),
            .I(N__30743));
    LocalMux I__5463 (
            .O(N__30752),
            .I(N__30743));
    InMux I__5462 (
            .O(N__30751),
            .I(N__30740));
    Odrv4 I__5461 (
            .O(N__30748),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__5460 (
            .O(N__30743),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__5459 (
            .O(N__30740),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__5458 (
            .O(N__30733),
            .I(N__30730));
    LocalMux I__5457 (
            .O(N__30730),
            .I(N__30725));
    InMux I__5456 (
            .O(N__30729),
            .I(N__30720));
    InMux I__5455 (
            .O(N__30728),
            .I(N__30720));
    Span4Mux_v I__5454 (
            .O(N__30725),
            .I(N__30717));
    LocalMux I__5453 (
            .O(N__30720),
            .I(N__30714));
    Odrv4 I__5452 (
            .O(N__30717),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__5451 (
            .O(N__30714),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__5450 (
            .O(N__30709),
            .I(N__30706));
    InMux I__5449 (
            .O(N__30706),
            .I(N__30703));
    LocalMux I__5448 (
            .O(N__30703),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    CascadeMux I__5447 (
            .O(N__30700),
            .I(N__30697));
    InMux I__5446 (
            .O(N__30697),
            .I(N__30691));
    InMux I__5445 (
            .O(N__30696),
            .I(N__30691));
    LocalMux I__5444 (
            .O(N__30691),
            .I(N__30688));
    Span4Mux_h I__5443 (
            .O(N__30688),
            .I(N__30685));
    Odrv4 I__5442 (
            .O(N__30685),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__5441 (
            .O(N__30682),
            .I(N__30679));
    LocalMux I__5440 (
            .O(N__30679),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    InMux I__5439 (
            .O(N__30676),
            .I(N__30673));
    LocalMux I__5438 (
            .O(N__30673),
            .I(N__30670));
    Span4Mux_h I__5437 (
            .O(N__30670),
            .I(N__30665));
    InMux I__5436 (
            .O(N__30669),
            .I(N__30660));
    InMux I__5435 (
            .O(N__30668),
            .I(N__30660));
    Span4Mux_v I__5434 (
            .O(N__30665),
            .I(N__30654));
    LocalMux I__5433 (
            .O(N__30660),
            .I(N__30654));
    InMux I__5432 (
            .O(N__30659),
            .I(N__30651));
    Odrv4 I__5431 (
            .O(N__30654),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5430 (
            .O(N__30651),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5429 (
            .O(N__30646),
            .I(N__30643));
    LocalMux I__5428 (
            .O(N__30643),
            .I(N__30640));
    Span4Mux_v I__5427 (
            .O(N__30640),
            .I(N__30636));
    InMux I__5426 (
            .O(N__30639),
            .I(N__30633));
    Odrv4 I__5425 (
            .O(N__30636),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__5424 (
            .O(N__30633),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__5423 (
            .O(N__30628),
            .I(N__30622));
    InMux I__5422 (
            .O(N__30627),
            .I(N__30622));
    LocalMux I__5421 (
            .O(N__30622),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__5420 (
            .O(N__30619),
            .I(N__30614));
    InMux I__5419 (
            .O(N__30618),
            .I(N__30608));
    InMux I__5418 (
            .O(N__30617),
            .I(N__30608));
    LocalMux I__5417 (
            .O(N__30614),
            .I(N__30605));
    InMux I__5416 (
            .O(N__30613),
            .I(N__30602));
    LocalMux I__5415 (
            .O(N__30608),
            .I(N__30599));
    Span4Mux_v I__5414 (
            .O(N__30605),
            .I(N__30596));
    LocalMux I__5413 (
            .O(N__30602),
            .I(N__30593));
    Span4Mux_h I__5412 (
            .O(N__30599),
            .I(N__30590));
    Span4Mux_h I__5411 (
            .O(N__30596),
            .I(N__30585));
    Span4Mux_h I__5410 (
            .O(N__30593),
            .I(N__30585));
    Odrv4 I__5409 (
            .O(N__30590),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__5408 (
            .O(N__30585),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__5407 (
            .O(N__30580),
            .I(N__30577));
    LocalMux I__5406 (
            .O(N__30577),
            .I(N__30574));
    Span4Mux_v I__5405 (
            .O(N__30574),
            .I(N__30570));
    InMux I__5404 (
            .O(N__30573),
            .I(N__30567));
    Odrv4 I__5403 (
            .O(N__30570),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__5402 (
            .O(N__30567),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    InMux I__5401 (
            .O(N__30562),
            .I(N__30543));
    InMux I__5400 (
            .O(N__30561),
            .I(N__30543));
    InMux I__5399 (
            .O(N__30560),
            .I(N__30538));
    InMux I__5398 (
            .O(N__30559),
            .I(N__30538));
    CascadeMux I__5397 (
            .O(N__30558),
            .I(N__30531));
    InMux I__5396 (
            .O(N__30557),
            .I(N__30523));
    InMux I__5395 (
            .O(N__30556),
            .I(N__30516));
    InMux I__5394 (
            .O(N__30555),
            .I(N__30516));
    InMux I__5393 (
            .O(N__30554),
            .I(N__30516));
    InMux I__5392 (
            .O(N__30553),
            .I(N__30505));
    InMux I__5391 (
            .O(N__30552),
            .I(N__30505));
    InMux I__5390 (
            .O(N__30551),
            .I(N__30505));
    InMux I__5389 (
            .O(N__30550),
            .I(N__30505));
    InMux I__5388 (
            .O(N__30549),
            .I(N__30505));
    CascadeMux I__5387 (
            .O(N__30548),
            .I(N__30494));
    LocalMux I__5386 (
            .O(N__30543),
            .I(N__30487));
    LocalMux I__5385 (
            .O(N__30538),
            .I(N__30484));
    InMux I__5384 (
            .O(N__30537),
            .I(N__30467));
    InMux I__5383 (
            .O(N__30536),
            .I(N__30467));
    InMux I__5382 (
            .O(N__30535),
            .I(N__30467));
    InMux I__5381 (
            .O(N__30534),
            .I(N__30467));
    InMux I__5380 (
            .O(N__30531),
            .I(N__30467));
    InMux I__5379 (
            .O(N__30530),
            .I(N__30467));
    InMux I__5378 (
            .O(N__30529),
            .I(N__30467));
    InMux I__5377 (
            .O(N__30528),
            .I(N__30467));
    InMux I__5376 (
            .O(N__30527),
            .I(N__30462));
    InMux I__5375 (
            .O(N__30526),
            .I(N__30462));
    LocalMux I__5374 (
            .O(N__30523),
            .I(N__30455));
    LocalMux I__5373 (
            .O(N__30516),
            .I(N__30455));
    LocalMux I__5372 (
            .O(N__30505),
            .I(N__30455));
    InMux I__5371 (
            .O(N__30504),
            .I(N__30442));
    InMux I__5370 (
            .O(N__30503),
            .I(N__30442));
    InMux I__5369 (
            .O(N__30502),
            .I(N__30442));
    InMux I__5368 (
            .O(N__30501),
            .I(N__30442));
    InMux I__5367 (
            .O(N__30500),
            .I(N__30442));
    InMux I__5366 (
            .O(N__30499),
            .I(N__30442));
    InMux I__5365 (
            .O(N__30498),
            .I(N__30416));
    InMux I__5364 (
            .O(N__30497),
            .I(N__30409));
    InMux I__5363 (
            .O(N__30494),
            .I(N__30409));
    InMux I__5362 (
            .O(N__30493),
            .I(N__30409));
    InMux I__5361 (
            .O(N__30492),
            .I(N__30402));
    InMux I__5360 (
            .O(N__30491),
            .I(N__30402));
    InMux I__5359 (
            .O(N__30490),
            .I(N__30402));
    Span4Mux_v I__5358 (
            .O(N__30487),
            .I(N__30389));
    Span4Mux_v I__5357 (
            .O(N__30484),
            .I(N__30389));
    LocalMux I__5356 (
            .O(N__30467),
            .I(N__30389));
    LocalMux I__5355 (
            .O(N__30462),
            .I(N__30389));
    Span4Mux_v I__5354 (
            .O(N__30455),
            .I(N__30389));
    LocalMux I__5353 (
            .O(N__30442),
            .I(N__30389));
    InMux I__5352 (
            .O(N__30441),
            .I(N__30378));
    InMux I__5351 (
            .O(N__30440),
            .I(N__30378));
    InMux I__5350 (
            .O(N__30439),
            .I(N__30378));
    InMux I__5349 (
            .O(N__30438),
            .I(N__30378));
    InMux I__5348 (
            .O(N__30437),
            .I(N__30378));
    InMux I__5347 (
            .O(N__30436),
            .I(N__30369));
    InMux I__5346 (
            .O(N__30435),
            .I(N__30369));
    InMux I__5345 (
            .O(N__30434),
            .I(N__30369));
    InMux I__5344 (
            .O(N__30433),
            .I(N__30369));
    InMux I__5343 (
            .O(N__30432),
            .I(N__30365));
    InMux I__5342 (
            .O(N__30431),
            .I(N__30358));
    InMux I__5341 (
            .O(N__30430),
            .I(N__30358));
    InMux I__5340 (
            .O(N__30429),
            .I(N__30358));
    InMux I__5339 (
            .O(N__30428),
            .I(N__30347));
    InMux I__5338 (
            .O(N__30427),
            .I(N__30347));
    InMux I__5337 (
            .O(N__30426),
            .I(N__30347));
    InMux I__5336 (
            .O(N__30425),
            .I(N__30347));
    InMux I__5335 (
            .O(N__30424),
            .I(N__30343));
    InMux I__5334 (
            .O(N__30423),
            .I(N__30336));
    InMux I__5333 (
            .O(N__30422),
            .I(N__30336));
    InMux I__5332 (
            .O(N__30421),
            .I(N__30336));
    InMux I__5331 (
            .O(N__30420),
            .I(N__30331));
    InMux I__5330 (
            .O(N__30419),
            .I(N__30331));
    LocalMux I__5329 (
            .O(N__30416),
            .I(N__30306));
    LocalMux I__5328 (
            .O(N__30409),
            .I(N__30306));
    LocalMux I__5327 (
            .O(N__30402),
            .I(N__30306));
    Span4Mux_h I__5326 (
            .O(N__30389),
            .I(N__30306));
    LocalMux I__5325 (
            .O(N__30378),
            .I(N__30306));
    LocalMux I__5324 (
            .O(N__30369),
            .I(N__30306));
    InMux I__5323 (
            .O(N__30368),
            .I(N__30299));
    LocalMux I__5322 (
            .O(N__30365),
            .I(N__30296));
    LocalMux I__5321 (
            .O(N__30358),
            .I(N__30293));
    InMux I__5320 (
            .O(N__30357),
            .I(N__30288));
    InMux I__5319 (
            .O(N__30356),
            .I(N__30288));
    LocalMux I__5318 (
            .O(N__30347),
            .I(N__30285));
    InMux I__5317 (
            .O(N__30346),
            .I(N__30282));
    LocalMux I__5316 (
            .O(N__30343),
            .I(N__30275));
    LocalMux I__5315 (
            .O(N__30336),
            .I(N__30275));
    LocalMux I__5314 (
            .O(N__30331),
            .I(N__30275));
    InMux I__5313 (
            .O(N__30330),
            .I(N__30270));
    InMux I__5312 (
            .O(N__30329),
            .I(N__30270));
    InMux I__5311 (
            .O(N__30328),
            .I(N__30267));
    InMux I__5310 (
            .O(N__30327),
            .I(N__30260));
    InMux I__5309 (
            .O(N__30326),
            .I(N__30260));
    InMux I__5308 (
            .O(N__30325),
            .I(N__30260));
    InMux I__5307 (
            .O(N__30324),
            .I(N__30255));
    InMux I__5306 (
            .O(N__30323),
            .I(N__30255));
    InMux I__5305 (
            .O(N__30322),
            .I(N__30248));
    InMux I__5304 (
            .O(N__30321),
            .I(N__30248));
    InMux I__5303 (
            .O(N__30320),
            .I(N__30248));
    InMux I__5302 (
            .O(N__30319),
            .I(N__30238));
    Span4Mux_v I__5301 (
            .O(N__30306),
            .I(N__30235));
    InMux I__5300 (
            .O(N__30305),
            .I(N__30228));
    InMux I__5299 (
            .O(N__30304),
            .I(N__30228));
    InMux I__5298 (
            .O(N__30303),
            .I(N__30228));
    InMux I__5297 (
            .O(N__30302),
            .I(N__30222));
    LocalMux I__5296 (
            .O(N__30299),
            .I(N__30210));
    Span4Mux_v I__5295 (
            .O(N__30296),
            .I(N__30210));
    Span4Mux_v I__5294 (
            .O(N__30293),
            .I(N__30210));
    LocalMux I__5293 (
            .O(N__30288),
            .I(N__30210));
    Span4Mux_v I__5292 (
            .O(N__30285),
            .I(N__30205));
    LocalMux I__5291 (
            .O(N__30282),
            .I(N__30205));
    Span4Mux_h I__5290 (
            .O(N__30275),
            .I(N__30198));
    LocalMux I__5289 (
            .O(N__30270),
            .I(N__30198));
    LocalMux I__5288 (
            .O(N__30267),
            .I(N__30198));
    LocalMux I__5287 (
            .O(N__30260),
            .I(N__30191));
    LocalMux I__5286 (
            .O(N__30255),
            .I(N__30191));
    LocalMux I__5285 (
            .O(N__30248),
            .I(N__30191));
    InMux I__5284 (
            .O(N__30247),
            .I(N__30188));
    InMux I__5283 (
            .O(N__30246),
            .I(N__30183));
    InMux I__5282 (
            .O(N__30245),
            .I(N__30183));
    InMux I__5281 (
            .O(N__30244),
            .I(N__30180));
    InMux I__5280 (
            .O(N__30243),
            .I(N__30177));
    InMux I__5279 (
            .O(N__30242),
            .I(N__30172));
    InMux I__5278 (
            .O(N__30241),
            .I(N__30172));
    LocalMux I__5277 (
            .O(N__30238),
            .I(N__30165));
    Sp12to4 I__5276 (
            .O(N__30235),
            .I(N__30165));
    LocalMux I__5275 (
            .O(N__30228),
            .I(N__30165));
    InMux I__5274 (
            .O(N__30227),
            .I(N__30160));
    InMux I__5273 (
            .O(N__30226),
            .I(N__30160));
    InMux I__5272 (
            .O(N__30225),
            .I(N__30157));
    LocalMux I__5271 (
            .O(N__30222),
            .I(N__30154));
    InMux I__5270 (
            .O(N__30221),
            .I(N__30147));
    InMux I__5269 (
            .O(N__30220),
            .I(N__30147));
    InMux I__5268 (
            .O(N__30219),
            .I(N__30147));
    Span4Mux_h I__5267 (
            .O(N__30210),
            .I(N__30142));
    Span4Mux_h I__5266 (
            .O(N__30205),
            .I(N__30142));
    Span4Mux_h I__5265 (
            .O(N__30198),
            .I(N__30139));
    Span12Mux_v I__5264 (
            .O(N__30191),
            .I(N__30136));
    LocalMux I__5263 (
            .O(N__30188),
            .I(N__30123));
    LocalMux I__5262 (
            .O(N__30183),
            .I(N__30123));
    LocalMux I__5261 (
            .O(N__30180),
            .I(N__30123));
    LocalMux I__5260 (
            .O(N__30177),
            .I(N__30123));
    LocalMux I__5259 (
            .O(N__30172),
            .I(N__30123));
    Span12Mux_h I__5258 (
            .O(N__30165),
            .I(N__30123));
    LocalMux I__5257 (
            .O(N__30160),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5256 (
            .O(N__30157),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5255 (
            .O(N__30154),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5254 (
            .O(N__30147),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5253 (
            .O(N__30142),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5252 (
            .O(N__30139),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__5251 (
            .O(N__30136),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__5250 (
            .O(N__30123),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    CEMux I__5249 (
            .O(N__30106),
            .I(N__30073));
    CEMux I__5248 (
            .O(N__30105),
            .I(N__30073));
    CEMux I__5247 (
            .O(N__30104),
            .I(N__30073));
    CEMux I__5246 (
            .O(N__30103),
            .I(N__30073));
    CEMux I__5245 (
            .O(N__30102),
            .I(N__30073));
    CEMux I__5244 (
            .O(N__30101),
            .I(N__30073));
    CEMux I__5243 (
            .O(N__30100),
            .I(N__30073));
    CEMux I__5242 (
            .O(N__30099),
            .I(N__30073));
    CEMux I__5241 (
            .O(N__30098),
            .I(N__30073));
    CEMux I__5240 (
            .O(N__30097),
            .I(N__30073));
    CEMux I__5239 (
            .O(N__30096),
            .I(N__30073));
    GlobalMux I__5238 (
            .O(N__30073),
            .I(N__30070));
    gio2CtrlBuf I__5237 (
            .O(N__30070),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__5236 (
            .O(N__30067),
            .I(N__30064));
    LocalMux I__5235 (
            .O(N__30064),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    CascadeMux I__5234 (
            .O(N__30061),
            .I(N__30058));
    InMux I__5233 (
            .O(N__30058),
            .I(N__30052));
    InMux I__5232 (
            .O(N__30057),
            .I(N__30052));
    LocalMux I__5231 (
            .O(N__30052),
            .I(N__30049));
    Span4Mux_v I__5230 (
            .O(N__30049),
            .I(N__30046));
    Odrv4 I__5229 (
            .O(N__30046),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__5228 (
            .O(N__30043),
            .I(N__30037));
    InMux I__5227 (
            .O(N__30042),
            .I(N__30037));
    LocalMux I__5226 (
            .O(N__30037),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__5225 (
            .O(N__30034),
            .I(N__30031));
    InMux I__5224 (
            .O(N__30031),
            .I(N__30028));
    LocalMux I__5223 (
            .O(N__30028),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    InMux I__5222 (
            .O(N__30025),
            .I(N__30022));
    LocalMux I__5221 (
            .O(N__30022),
            .I(N__30018));
    InMux I__5220 (
            .O(N__30021),
            .I(N__30015));
    Span4Mux_h I__5219 (
            .O(N__30018),
            .I(N__30010));
    LocalMux I__5218 (
            .O(N__30015),
            .I(N__30010));
    Odrv4 I__5217 (
            .O(N__30010),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__5216 (
            .O(N__30007),
            .I(N__30003));
    InMux I__5215 (
            .O(N__30006),
            .I(N__30000));
    InMux I__5214 (
            .O(N__30003),
            .I(N__29997));
    LocalMux I__5213 (
            .O(N__30000),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    LocalMux I__5212 (
            .O(N__29997),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__5211 (
            .O(N__29992),
            .I(N__29989));
    InMux I__5210 (
            .O(N__29989),
            .I(N__29986));
    LocalMux I__5209 (
            .O(N__29986),
            .I(N__29983));
    Odrv4 I__5208 (
            .O(N__29983),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__5207 (
            .O(N__29980),
            .I(N__29976));
    InMux I__5206 (
            .O(N__29979),
            .I(N__29973));
    LocalMux I__5205 (
            .O(N__29976),
            .I(N__29970));
    LocalMux I__5204 (
            .O(N__29973),
            .I(N__29967));
    Span4Mux_v I__5203 (
            .O(N__29970),
            .I(N__29964));
    Span12Mux_v I__5202 (
            .O(N__29967),
            .I(N__29961));
    Span4Mux_h I__5201 (
            .O(N__29964),
            .I(N__29958));
    Odrv12 I__5200 (
            .O(N__29961),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__5199 (
            .O(N__29958),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5198 (
            .O(N__29953),
            .I(N__29950));
    LocalMux I__5197 (
            .O(N__29950),
            .I(N__29946));
    InMux I__5196 (
            .O(N__29949),
            .I(N__29943));
    Span4Mux_h I__5195 (
            .O(N__29946),
            .I(N__29940));
    LocalMux I__5194 (
            .O(N__29943),
            .I(N__29937));
    Span4Mux_h I__5193 (
            .O(N__29940),
            .I(N__29934));
    Span12Mux_s7_h I__5192 (
            .O(N__29937),
            .I(N__29931));
    Odrv4 I__5191 (
            .O(N__29934),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv12 I__5190 (
            .O(N__29931),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__5189 (
            .O(N__29926),
            .I(N__29922));
    InMux I__5188 (
            .O(N__29925),
            .I(N__29919));
    LocalMux I__5187 (
            .O(N__29922),
            .I(N__29916));
    LocalMux I__5186 (
            .O(N__29919),
            .I(N__29913));
    Span4Mux_h I__5185 (
            .O(N__29916),
            .I(N__29910));
    Span4Mux_v I__5184 (
            .O(N__29913),
            .I(N__29907));
    Sp12to4 I__5183 (
            .O(N__29910),
            .I(N__29904));
    Sp12to4 I__5182 (
            .O(N__29907),
            .I(N__29899));
    Span12Mux_v I__5181 (
            .O(N__29904),
            .I(N__29899));
    Odrv12 I__5180 (
            .O(N__29899),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__5179 (
            .O(N__29896),
            .I(N__29893));
    LocalMux I__5178 (
            .O(N__29893),
            .I(N__29890));
    Odrv12 I__5177 (
            .O(N__29890),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__5176 (
            .O(N__29887),
            .I(N__29884));
    InMux I__5175 (
            .O(N__29884),
            .I(N__29881));
    LocalMux I__5174 (
            .O(N__29881),
            .I(N__29878));
    Odrv12 I__5173 (
            .O(N__29878),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__5172 (
            .O(N__29875),
            .I(N__29872));
    LocalMux I__5171 (
            .O(N__29872),
            .I(N__29869));
    Odrv4 I__5170 (
            .O(N__29869),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    CascadeMux I__5169 (
            .O(N__29866),
            .I(N__29863));
    InMux I__5168 (
            .O(N__29863),
            .I(N__29860));
    LocalMux I__5167 (
            .O(N__29860),
            .I(N__29857));
    Odrv4 I__5166 (
            .O(N__29857),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    InMux I__5165 (
            .O(N__29854),
            .I(N__29851));
    LocalMux I__5164 (
            .O(N__29851),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    CascadeMux I__5163 (
            .O(N__29848),
            .I(N__29845));
    InMux I__5162 (
            .O(N__29845),
            .I(N__29842));
    LocalMux I__5161 (
            .O(N__29842),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__5160 (
            .O(N__29839),
            .I(N__29836));
    LocalMux I__5159 (
            .O(N__29836),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    InMux I__5158 (
            .O(N__29833),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__5157 (
            .O(N__29830),
            .I(N__29827));
    InMux I__5156 (
            .O(N__29827),
            .I(N__29824));
    LocalMux I__5155 (
            .O(N__29824),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    CascadeMux I__5154 (
            .O(N__29821),
            .I(N__29818));
    InMux I__5153 (
            .O(N__29818),
            .I(N__29815));
    LocalMux I__5152 (
            .O(N__29815),
            .I(N__29812));
    Odrv12 I__5151 (
            .O(N__29812),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__5150 (
            .O(N__29809),
            .I(N__29806));
    LocalMux I__5149 (
            .O(N__29806),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__5148 (
            .O(N__29803),
            .I(N__29800));
    InMux I__5147 (
            .O(N__29800),
            .I(N__29797));
    LocalMux I__5146 (
            .O(N__29797),
            .I(N__29794));
    Odrv4 I__5145 (
            .O(N__29794),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__5144 (
            .O(N__29791),
            .I(N__29788));
    LocalMux I__5143 (
            .O(N__29788),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__5142 (
            .O(N__29785),
            .I(N__29782));
    LocalMux I__5141 (
            .O(N__29782),
            .I(N__29779));
    Odrv4 I__5140 (
            .O(N__29779),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__5139 (
            .O(N__29776),
            .I(N__29773));
    InMux I__5138 (
            .O(N__29773),
            .I(N__29770));
    LocalMux I__5137 (
            .O(N__29770),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__5136 (
            .O(N__29767),
            .I(N__29764));
    LocalMux I__5135 (
            .O(N__29764),
            .I(N__29761));
    Span4Mux_v I__5134 (
            .O(N__29761),
            .I(N__29758));
    Span4Mux_h I__5133 (
            .O(N__29758),
            .I(N__29755));
    Odrv4 I__5132 (
            .O(N__29755),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__5131 (
            .O(N__29752),
            .I(N__29749));
    InMux I__5130 (
            .O(N__29749),
            .I(N__29746));
    LocalMux I__5129 (
            .O(N__29746),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__5128 (
            .O(N__29743),
            .I(N__29740));
    LocalMux I__5127 (
            .O(N__29740),
            .I(N__29737));
    Odrv4 I__5126 (
            .O(N__29737),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__5125 (
            .O(N__29734),
            .I(N__29731));
    InMux I__5124 (
            .O(N__29731),
            .I(N__29728));
    LocalMux I__5123 (
            .O(N__29728),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__5122 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__5121 (
            .O(N__29722),
            .I(N__29719));
    Odrv4 I__5120 (
            .O(N__29719),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__5119 (
            .O(N__29716),
            .I(N__29713));
    InMux I__5118 (
            .O(N__29713),
            .I(N__29710));
    LocalMux I__5117 (
            .O(N__29710),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__5116 (
            .O(N__29707),
            .I(N__29704));
    LocalMux I__5115 (
            .O(N__29704),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    CascadeMux I__5114 (
            .O(N__29701),
            .I(N__29698));
    InMux I__5113 (
            .O(N__29698),
            .I(N__29695));
    LocalMux I__5112 (
            .O(N__29695),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__5111 (
            .O(N__29692),
            .I(N__29689));
    LocalMux I__5110 (
            .O(N__29689),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__5109 (
            .O(N__29686),
            .I(N__29683));
    InMux I__5108 (
            .O(N__29683),
            .I(N__29680));
    LocalMux I__5107 (
            .O(N__29680),
            .I(N__29677));
    Odrv4 I__5106 (
            .O(N__29677),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__5105 (
            .O(N__29674),
            .I(N__29671));
    LocalMux I__5104 (
            .O(N__29671),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__5103 (
            .O(N__29668),
            .I(N__29665));
    InMux I__5102 (
            .O(N__29665),
            .I(N__29662));
    LocalMux I__5101 (
            .O(N__29662),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__5100 (
            .O(N__29659),
            .I(N__29656));
    LocalMux I__5099 (
            .O(N__29656),
            .I(N__29653));
    Span4Mux_h I__5098 (
            .O(N__29653),
            .I(N__29650));
    Odrv4 I__5097 (
            .O(N__29650),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__5096 (
            .O(N__29647),
            .I(N__29644));
    InMux I__5095 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__5094 (
            .O(N__29641),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__5093 (
            .O(N__29638),
            .I(N__29635));
    LocalMux I__5092 (
            .O(N__29635),
            .I(N__29632));
    Odrv12 I__5091 (
            .O(N__29632),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__5090 (
            .O(N__29629),
            .I(N__29626));
    InMux I__5089 (
            .O(N__29626),
            .I(N__29623));
    LocalMux I__5088 (
            .O(N__29623),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__5087 (
            .O(N__29620),
            .I(N__29617));
    LocalMux I__5086 (
            .O(N__29617),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__5085 (
            .O(N__29614),
            .I(N__29611));
    InMux I__5084 (
            .O(N__29611),
            .I(N__29608));
    LocalMux I__5083 (
            .O(N__29608),
            .I(N__29605));
    Odrv4 I__5082 (
            .O(N__29605),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__5081 (
            .O(N__29602),
            .I(N__29599));
    InMux I__5080 (
            .O(N__29599),
            .I(N__29596));
    LocalMux I__5079 (
            .O(N__29596),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    InMux I__5078 (
            .O(N__29593),
            .I(N__29590));
    LocalMux I__5077 (
            .O(N__29590),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__5076 (
            .O(N__29587),
            .I(N__29584));
    InMux I__5075 (
            .O(N__29584),
            .I(N__29581));
    LocalMux I__5074 (
            .O(N__29581),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__5073 (
            .O(N__29578),
            .I(N__29575));
    LocalMux I__5072 (
            .O(N__29575),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__5071 (
            .O(N__29572),
            .I(N__29569));
    InMux I__5070 (
            .O(N__29569),
            .I(N__29566));
    LocalMux I__5069 (
            .O(N__29566),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    InMux I__5068 (
            .O(N__29563),
            .I(N__29560));
    LocalMux I__5067 (
            .O(N__29560),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__5066 (
            .O(N__29557),
            .I(N__29554));
    LocalMux I__5065 (
            .O(N__29554),
            .I(N__29551));
    Odrv4 I__5064 (
            .O(N__29551),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__5063 (
            .O(N__29548),
            .I(N__29545));
    InMux I__5062 (
            .O(N__29545),
            .I(N__29542));
    LocalMux I__5061 (
            .O(N__29542),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__5060 (
            .O(N__29539),
            .I(N__29534));
    InMux I__5059 (
            .O(N__29538),
            .I(N__29531));
    InMux I__5058 (
            .O(N__29537),
            .I(N__29528));
    LocalMux I__5057 (
            .O(N__29534),
            .I(N__29523));
    LocalMux I__5056 (
            .O(N__29531),
            .I(N__29523));
    LocalMux I__5055 (
            .O(N__29528),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__5054 (
            .O(N__29523),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__5053 (
            .O(N__29518),
            .I(N__29514));
    InMux I__5052 (
            .O(N__29517),
            .I(N__29511));
    LocalMux I__5051 (
            .O(N__29514),
            .I(N__29508));
    LocalMux I__5050 (
            .O(N__29511),
            .I(N__29504));
    Span4Mux_v I__5049 (
            .O(N__29508),
            .I(N__29501));
    InMux I__5048 (
            .O(N__29507),
            .I(N__29498));
    Span4Mux_h I__5047 (
            .O(N__29504),
            .I(N__29495));
    Sp12to4 I__5046 (
            .O(N__29501),
            .I(N__29489));
    LocalMux I__5045 (
            .O(N__29498),
            .I(N__29489));
    Span4Mux_h I__5044 (
            .O(N__29495),
            .I(N__29486));
    InMux I__5043 (
            .O(N__29494),
            .I(N__29483));
    Odrv12 I__5042 (
            .O(N__29489),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__5041 (
            .O(N__29486),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__5040 (
            .O(N__29483),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CascadeMux I__5039 (
            .O(N__29476),
            .I(N__29472));
    InMux I__5038 (
            .O(N__29475),
            .I(N__29467));
    InMux I__5037 (
            .O(N__29472),
            .I(N__29467));
    LocalMux I__5036 (
            .O(N__29467),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__5035 (
            .O(N__29464),
            .I(N__29459));
    InMux I__5034 (
            .O(N__29463),
            .I(N__29454));
    InMux I__5033 (
            .O(N__29462),
            .I(N__29454));
    LocalMux I__5032 (
            .O(N__29459),
            .I(N__29451));
    LocalMux I__5031 (
            .O(N__29454),
            .I(N__29448));
    Span4Mux_h I__5030 (
            .O(N__29451),
            .I(N__29442));
    Span4Mux_v I__5029 (
            .O(N__29448),
            .I(N__29442));
    InMux I__5028 (
            .O(N__29447),
            .I(N__29439));
    Odrv4 I__5027 (
            .O(N__29442),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__5026 (
            .O(N__29439),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__5025 (
            .O(N__29434),
            .I(N__29431));
    LocalMux I__5024 (
            .O(N__29431),
            .I(N__29427));
    InMux I__5023 (
            .O(N__29430),
            .I(N__29424));
    Odrv4 I__5022 (
            .O(N__29427),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__5021 (
            .O(N__29424),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__5020 (
            .O(N__29419),
            .I(N__29413));
    InMux I__5019 (
            .O(N__29418),
            .I(N__29413));
    LocalMux I__5018 (
            .O(N__29413),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__5017 (
            .O(N__29410),
            .I(N__29407));
    LocalMux I__5016 (
            .O(N__29407),
            .I(N__29403));
    InMux I__5015 (
            .O(N__29406),
            .I(N__29400));
    Odrv4 I__5014 (
            .O(N__29403),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    LocalMux I__5013 (
            .O(N__29400),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__5012 (
            .O(N__29395),
            .I(N__29390));
    InMux I__5011 (
            .O(N__29394),
            .I(N__29385));
    InMux I__5010 (
            .O(N__29393),
            .I(N__29385));
    LocalMux I__5009 (
            .O(N__29390),
            .I(N__29379));
    LocalMux I__5008 (
            .O(N__29385),
            .I(N__29379));
    InMux I__5007 (
            .O(N__29384),
            .I(N__29376));
    Span4Mux_v I__5006 (
            .O(N__29379),
            .I(N__29371));
    LocalMux I__5005 (
            .O(N__29376),
            .I(N__29371));
    Span4Mux_h I__5004 (
            .O(N__29371),
            .I(N__29368));
    Odrv4 I__5003 (
            .O(N__29368),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    CascadeMux I__5002 (
            .O(N__29365),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    InMux I__5001 (
            .O(N__29362),
            .I(N__29357));
    InMux I__5000 (
            .O(N__29361),
            .I(N__29352));
    InMux I__4999 (
            .O(N__29360),
            .I(N__29352));
    LocalMux I__4998 (
            .O(N__29357),
            .I(N__29346));
    LocalMux I__4997 (
            .O(N__29352),
            .I(N__29346));
    InMux I__4996 (
            .O(N__29351),
            .I(N__29343));
    Span4Mux_v I__4995 (
            .O(N__29346),
            .I(N__29338));
    LocalMux I__4994 (
            .O(N__29343),
            .I(N__29338));
    Span4Mux_h I__4993 (
            .O(N__29338),
            .I(N__29335));
    Odrv4 I__4992 (
            .O(N__29335),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__4991 (
            .O(N__29332),
            .I(N__29328));
    InMux I__4990 (
            .O(N__29331),
            .I(N__29325));
    LocalMux I__4989 (
            .O(N__29328),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__4988 (
            .O(N__29325),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    CascadeMux I__4987 (
            .O(N__29320),
            .I(N__29317));
    InMux I__4986 (
            .O(N__29317),
            .I(N__29314));
    LocalMux I__4985 (
            .O(N__29314),
            .I(N__29311));
    Odrv12 I__4984 (
            .O(N__29311),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    InMux I__4983 (
            .O(N__29308),
            .I(N__29305));
    LocalMux I__4982 (
            .O(N__29305),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__4981 (
            .O(N__29302),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_));
    InMux I__4980 (
            .O(N__29299),
            .I(N__29296));
    LocalMux I__4979 (
            .O(N__29296),
            .I(N__29293));
    Odrv4 I__4978 (
            .O(N__29293),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__4977 (
            .O(N__29290),
            .I(N__29287));
    InMux I__4976 (
            .O(N__29287),
            .I(N__29284));
    LocalMux I__4975 (
            .O(N__29284),
            .I(N__29281));
    Span4Mux_h I__4974 (
            .O(N__29281),
            .I(N__29278));
    Odrv4 I__4973 (
            .O(N__29278),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CEMux I__4972 (
            .O(N__29275),
            .I(N__29271));
    CEMux I__4971 (
            .O(N__29274),
            .I(N__29268));
    LocalMux I__4970 (
            .O(N__29271),
            .I(N__29260));
    LocalMux I__4969 (
            .O(N__29268),
            .I(N__29260));
    CEMux I__4968 (
            .O(N__29267),
            .I(N__29257));
    CEMux I__4967 (
            .O(N__29266),
            .I(N__29249));
    CEMux I__4966 (
            .O(N__29265),
            .I(N__29243));
    Span4Mux_v I__4965 (
            .O(N__29260),
            .I(N__29230));
    LocalMux I__4964 (
            .O(N__29257),
            .I(N__29230));
    CEMux I__4963 (
            .O(N__29256),
            .I(N__29227));
    CEMux I__4962 (
            .O(N__29255),
            .I(N__29220));
    CEMux I__4961 (
            .O(N__29254),
            .I(N__29216));
    CEMux I__4960 (
            .O(N__29253),
            .I(N__29212));
    CEMux I__4959 (
            .O(N__29252),
            .I(N__29209));
    LocalMux I__4958 (
            .O(N__29249),
            .I(N__29206));
    CEMux I__4957 (
            .O(N__29248),
            .I(N__29203));
    CEMux I__4956 (
            .O(N__29247),
            .I(N__29200));
    CEMux I__4955 (
            .O(N__29246),
            .I(N__29197));
    LocalMux I__4954 (
            .O(N__29243),
            .I(N__29183));
    InMux I__4953 (
            .O(N__29242),
            .I(N__29174));
    InMux I__4952 (
            .O(N__29241),
            .I(N__29174));
    InMux I__4951 (
            .O(N__29240),
            .I(N__29174));
    InMux I__4950 (
            .O(N__29239),
            .I(N__29174));
    InMux I__4949 (
            .O(N__29238),
            .I(N__29167));
    InMux I__4948 (
            .O(N__29237),
            .I(N__29167));
    InMux I__4947 (
            .O(N__29236),
            .I(N__29167));
    CEMux I__4946 (
            .O(N__29235),
            .I(N__29164));
    Span4Mux_v I__4945 (
            .O(N__29230),
            .I(N__29159));
    LocalMux I__4944 (
            .O(N__29227),
            .I(N__29159));
    InMux I__4943 (
            .O(N__29226),
            .I(N__29150));
    InMux I__4942 (
            .O(N__29225),
            .I(N__29150));
    InMux I__4941 (
            .O(N__29224),
            .I(N__29150));
    InMux I__4940 (
            .O(N__29223),
            .I(N__29150));
    LocalMux I__4939 (
            .O(N__29220),
            .I(N__29146));
    CEMux I__4938 (
            .O(N__29219),
            .I(N__29143));
    LocalMux I__4937 (
            .O(N__29216),
            .I(N__29140));
    CEMux I__4936 (
            .O(N__29215),
            .I(N__29137));
    LocalMux I__4935 (
            .O(N__29212),
            .I(N__29132));
    LocalMux I__4934 (
            .O(N__29209),
            .I(N__29132));
    Span4Mux_h I__4933 (
            .O(N__29206),
            .I(N__29125));
    LocalMux I__4932 (
            .O(N__29203),
            .I(N__29125));
    LocalMux I__4931 (
            .O(N__29200),
            .I(N__29125));
    LocalMux I__4930 (
            .O(N__29197),
            .I(N__29114));
    InMux I__4929 (
            .O(N__29196),
            .I(N__29105));
    InMux I__4928 (
            .O(N__29195),
            .I(N__29105));
    InMux I__4927 (
            .O(N__29194),
            .I(N__29105));
    InMux I__4926 (
            .O(N__29193),
            .I(N__29105));
    InMux I__4925 (
            .O(N__29192),
            .I(N__29098));
    InMux I__4924 (
            .O(N__29191),
            .I(N__29098));
    InMux I__4923 (
            .O(N__29190),
            .I(N__29098));
    InMux I__4922 (
            .O(N__29189),
            .I(N__29089));
    InMux I__4921 (
            .O(N__29188),
            .I(N__29089));
    InMux I__4920 (
            .O(N__29187),
            .I(N__29089));
    InMux I__4919 (
            .O(N__29186),
            .I(N__29089));
    Span4Mux_h I__4918 (
            .O(N__29183),
            .I(N__29082));
    LocalMux I__4917 (
            .O(N__29174),
            .I(N__29082));
    LocalMux I__4916 (
            .O(N__29167),
            .I(N__29082));
    LocalMux I__4915 (
            .O(N__29164),
            .I(N__29077));
    Span4Mux_v I__4914 (
            .O(N__29159),
            .I(N__29077));
    LocalMux I__4913 (
            .O(N__29150),
            .I(N__29074));
    InMux I__4912 (
            .O(N__29149),
            .I(N__29071));
    Span4Mux_h I__4911 (
            .O(N__29146),
            .I(N__29068));
    LocalMux I__4910 (
            .O(N__29143),
            .I(N__29063));
    Span4Mux_v I__4909 (
            .O(N__29140),
            .I(N__29063));
    LocalMux I__4908 (
            .O(N__29137),
            .I(N__29058));
    Span4Mux_v I__4907 (
            .O(N__29132),
            .I(N__29058));
    Span4Mux_v I__4906 (
            .O(N__29125),
            .I(N__29055));
    InMux I__4905 (
            .O(N__29124),
            .I(N__29046));
    InMux I__4904 (
            .O(N__29123),
            .I(N__29046));
    InMux I__4903 (
            .O(N__29122),
            .I(N__29046));
    InMux I__4902 (
            .O(N__29121),
            .I(N__29046));
    InMux I__4901 (
            .O(N__29120),
            .I(N__29037));
    InMux I__4900 (
            .O(N__29119),
            .I(N__29037));
    InMux I__4899 (
            .O(N__29118),
            .I(N__29037));
    InMux I__4898 (
            .O(N__29117),
            .I(N__29037));
    Span4Mux_v I__4897 (
            .O(N__29114),
            .I(N__29034));
    LocalMux I__4896 (
            .O(N__29105),
            .I(N__29031));
    LocalMux I__4895 (
            .O(N__29098),
            .I(N__29020));
    LocalMux I__4894 (
            .O(N__29089),
            .I(N__29020));
    Span4Mux_v I__4893 (
            .O(N__29082),
            .I(N__29020));
    Span4Mux_h I__4892 (
            .O(N__29077),
            .I(N__29020));
    Span4Mux_v I__4891 (
            .O(N__29074),
            .I(N__29020));
    LocalMux I__4890 (
            .O(N__29071),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4889 (
            .O(N__29068),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4888 (
            .O(N__29063),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4887 (
            .O(N__29058),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4886 (
            .O(N__29055),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__4885 (
            .O(N__29046),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__4884 (
            .O(N__29037),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4883 (
            .O(N__29034),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4882 (
            .O(N__29031),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__4881 (
            .O(N__29020),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__4880 (
            .O(N__28999),
            .I(N__28996));
    LocalMux I__4879 (
            .O(N__28996),
            .I(N__28991));
    InMux I__4878 (
            .O(N__28995),
            .I(N__28988));
    InMux I__4877 (
            .O(N__28994),
            .I(N__28985));
    Span4Mux_v I__4876 (
            .O(N__28991),
            .I(N__28982));
    LocalMux I__4875 (
            .O(N__28988),
            .I(N__28979));
    LocalMux I__4874 (
            .O(N__28985),
            .I(N__28976));
    Span4Mux_h I__4873 (
            .O(N__28982),
            .I(N__28970));
    Span4Mux_h I__4872 (
            .O(N__28979),
            .I(N__28970));
    Span12Mux_h I__4871 (
            .O(N__28976),
            .I(N__28967));
    InMux I__4870 (
            .O(N__28975),
            .I(N__28964));
    Span4Mux_v I__4869 (
            .O(N__28970),
            .I(N__28961));
    Span12Mux_v I__4868 (
            .O(N__28967),
            .I(N__28958));
    LocalMux I__4867 (
            .O(N__28964),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__4866 (
            .O(N__28961),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__4865 (
            .O(N__28958),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__4864 (
            .O(N__28951),
            .I(N__28948));
    LocalMux I__4863 (
            .O(N__28948),
            .I(N__28942));
    InMux I__4862 (
            .O(N__28947),
            .I(N__28935));
    InMux I__4861 (
            .O(N__28946),
            .I(N__28935));
    InMux I__4860 (
            .O(N__28945),
            .I(N__28935));
    Span4Mux_v I__4859 (
            .O(N__28942),
            .I(N__28930));
    LocalMux I__4858 (
            .O(N__28935),
            .I(N__28930));
    Span4Mux_h I__4857 (
            .O(N__28930),
            .I(N__28927));
    Odrv4 I__4856 (
            .O(N__28927),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__4855 (
            .O(N__28924),
            .I(N__28921));
    LocalMux I__4854 (
            .O(N__28921),
            .I(N__28917));
    InMux I__4853 (
            .O(N__28920),
            .I(N__28914));
    Odrv4 I__4852 (
            .O(N__28917),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__4851 (
            .O(N__28914),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__4850 (
            .O(N__28909),
            .I(N__28904));
    InMux I__4849 (
            .O(N__28908),
            .I(N__28899));
    InMux I__4848 (
            .O(N__28907),
            .I(N__28899));
    LocalMux I__4847 (
            .O(N__28904),
            .I(N__28893));
    LocalMux I__4846 (
            .O(N__28899),
            .I(N__28893));
    InMux I__4845 (
            .O(N__28898),
            .I(N__28890));
    Span4Mux_v I__4844 (
            .O(N__28893),
            .I(N__28885));
    LocalMux I__4843 (
            .O(N__28890),
            .I(N__28885));
    Span4Mux_h I__4842 (
            .O(N__28885),
            .I(N__28882));
    Odrv4 I__4841 (
            .O(N__28882),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__4840 (
            .O(N__28879),
            .I(N__28875));
    InMux I__4839 (
            .O(N__28878),
            .I(N__28872));
    LocalMux I__4838 (
            .O(N__28875),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__4837 (
            .O(N__28872),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__4836 (
            .O(N__28867),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__4835 (
            .O(N__28864),
            .I(N__28860));
    CascadeMux I__4834 (
            .O(N__28863),
            .I(N__28857));
    LocalMux I__4833 (
            .O(N__28860),
            .I(N__28853));
    InMux I__4832 (
            .O(N__28857),
            .I(N__28850));
    InMux I__4831 (
            .O(N__28856),
            .I(N__28847));
    Span4Mux_h I__4830 (
            .O(N__28853),
            .I(N__28844));
    LocalMux I__4829 (
            .O(N__28850),
            .I(N__28841));
    LocalMux I__4828 (
            .O(N__28847),
            .I(N__28838));
    Span4Mux_v I__4827 (
            .O(N__28844),
            .I(N__28832));
    Span4Mux_h I__4826 (
            .O(N__28841),
            .I(N__28832));
    Span4Mux_h I__4825 (
            .O(N__28838),
            .I(N__28829));
    InMux I__4824 (
            .O(N__28837),
            .I(N__28826));
    Odrv4 I__4823 (
            .O(N__28832),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__4822 (
            .O(N__28829),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__4821 (
            .O(N__28826),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    CascadeMux I__4820 (
            .O(N__28819),
            .I(N__28815));
    InMux I__4819 (
            .O(N__28818),
            .I(N__28812));
    InMux I__4818 (
            .O(N__28815),
            .I(N__28809));
    LocalMux I__4817 (
            .O(N__28812),
            .I(N__28805));
    LocalMux I__4816 (
            .O(N__28809),
            .I(N__28802));
    InMux I__4815 (
            .O(N__28808),
            .I(N__28799));
    Span4Mux_v I__4814 (
            .O(N__28805),
            .I(N__28796));
    Odrv12 I__4813 (
            .O(N__28802),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__4812 (
            .O(N__28799),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__4811 (
            .O(N__28796),
            .I(\current_shift_inst.un4_control_input1_28 ));
    CascadeMux I__4810 (
            .O(N__28789),
            .I(N__28786));
    InMux I__4809 (
            .O(N__28786),
            .I(N__28783));
    LocalMux I__4808 (
            .O(N__28783),
            .I(N__28780));
    Odrv12 I__4807 (
            .O(N__28780),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__4806 (
            .O(N__28777),
            .I(N__28774));
    InMux I__4805 (
            .O(N__28774),
            .I(N__28771));
    LocalMux I__4804 (
            .O(N__28771),
            .I(N__28765));
    InMux I__4803 (
            .O(N__28770),
            .I(N__28762));
    InMux I__4802 (
            .O(N__28769),
            .I(N__28757));
    InMux I__4801 (
            .O(N__28768),
            .I(N__28757));
    Span4Mux_v I__4800 (
            .O(N__28765),
            .I(N__28754));
    LocalMux I__4799 (
            .O(N__28762),
            .I(N__28751));
    LocalMux I__4798 (
            .O(N__28757),
            .I(N__28748));
    Odrv4 I__4797 (
            .O(N__28754),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__4796 (
            .O(N__28751),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__4795 (
            .O(N__28748),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__4794 (
            .O(N__28741),
            .I(N__28737));
    CascadeMux I__4793 (
            .O(N__28740),
            .I(N__28734));
    LocalMux I__4792 (
            .O(N__28737),
            .I(N__28730));
    InMux I__4791 (
            .O(N__28734),
            .I(N__28727));
    InMux I__4790 (
            .O(N__28733),
            .I(N__28724));
    Span4Mux_v I__4789 (
            .O(N__28730),
            .I(N__28721));
    LocalMux I__4788 (
            .O(N__28727),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__4787 (
            .O(N__28724),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__4786 (
            .O(N__28721),
            .I(\current_shift_inst.un4_control_input1_30 ));
    CascadeMux I__4785 (
            .O(N__28714),
            .I(N__28711));
    InMux I__4784 (
            .O(N__28711),
            .I(N__28708));
    LocalMux I__4783 (
            .O(N__28708),
            .I(N__28705));
    Odrv12 I__4782 (
            .O(N__28705),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    IoInMux I__4781 (
            .O(N__28702),
            .I(N__28699));
    LocalMux I__4780 (
            .O(N__28699),
            .I(N__28696));
    IoSpan4Mux I__4779 (
            .O(N__28696),
            .I(N__28693));
    Span4Mux_s0_v I__4778 (
            .O(N__28693),
            .I(N__28690));
    Odrv4 I__4777 (
            .O(N__28690),
            .I(s3_phy_c));
    InMux I__4776 (
            .O(N__28687),
            .I(N__28684));
    LocalMux I__4775 (
            .O(N__28684),
            .I(N__28681));
    Glb2LocalMux I__4774 (
            .O(N__28681),
            .I(N__28678));
    GlobalMux I__4773 (
            .O(N__28678),
            .I(clk_12mhz));
    IoInMux I__4772 (
            .O(N__28675),
            .I(N__28672));
    LocalMux I__4771 (
            .O(N__28672),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__4770 (
            .O(N__28669),
            .I(N__28664));
    InMux I__4769 (
            .O(N__28668),
            .I(N__28661));
    InMux I__4768 (
            .O(N__28667),
            .I(N__28658));
    LocalMux I__4767 (
            .O(N__28664),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__4766 (
            .O(N__28661),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__4765 (
            .O(N__28658),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__4764 (
            .O(N__28651),
            .I(N__28647));
    InMux I__4763 (
            .O(N__28650),
            .I(N__28643));
    LocalMux I__4762 (
            .O(N__28647),
            .I(N__28640));
    InMux I__4761 (
            .O(N__28646),
            .I(N__28637));
    LocalMux I__4760 (
            .O(N__28643),
            .I(N__28633));
    Span4Mux_h I__4759 (
            .O(N__28640),
            .I(N__28628));
    LocalMux I__4758 (
            .O(N__28637),
            .I(N__28628));
    CascadeMux I__4757 (
            .O(N__28636),
            .I(N__28625));
    Span4Mux_h I__4756 (
            .O(N__28633),
            .I(N__28622));
    Span4Mux_h I__4755 (
            .O(N__28628),
            .I(N__28619));
    InMux I__4754 (
            .O(N__28625),
            .I(N__28616));
    Odrv4 I__4753 (
            .O(N__28622),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__4752 (
            .O(N__28619),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__4751 (
            .O(N__28616),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__4750 (
            .O(N__28609),
            .I(N__28606));
    LocalMux I__4749 (
            .O(N__28606),
            .I(N__28600));
    InMux I__4748 (
            .O(N__28605),
            .I(N__28595));
    InMux I__4747 (
            .O(N__28604),
            .I(N__28595));
    InMux I__4746 (
            .O(N__28603),
            .I(N__28592));
    Odrv4 I__4745 (
            .O(N__28600),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__4744 (
            .O(N__28595),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__4743 (
            .O(N__28592),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__4742 (
            .O(N__28585),
            .I(N__28581));
    CascadeMux I__4741 (
            .O(N__28584),
            .I(N__28578));
    InMux I__4740 (
            .O(N__28581),
            .I(N__28572));
    InMux I__4739 (
            .O(N__28578),
            .I(N__28569));
    InMux I__4738 (
            .O(N__28577),
            .I(N__28562));
    InMux I__4737 (
            .O(N__28576),
            .I(N__28562));
    InMux I__4736 (
            .O(N__28575),
            .I(N__28562));
    LocalMux I__4735 (
            .O(N__28572),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__4734 (
            .O(N__28569),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__4733 (
            .O(N__28562),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__4732 (
            .O(N__28555),
            .I(N__28551));
    InMux I__4731 (
            .O(N__28554),
            .I(N__28548));
    LocalMux I__4730 (
            .O(N__28551),
            .I(N__28542));
    LocalMux I__4729 (
            .O(N__28548),
            .I(N__28542));
    InMux I__4728 (
            .O(N__28547),
            .I(N__28539));
    Span4Mux_h I__4727 (
            .O(N__28542),
            .I(N__28536));
    LocalMux I__4726 (
            .O(N__28539),
            .I(N__28533));
    Odrv4 I__4725 (
            .O(N__28536),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv12 I__4724 (
            .O(N__28533),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__4723 (
            .O(N__28528),
            .I(N__28525));
    LocalMux I__4722 (
            .O(N__28525),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__4721 (
            .O(N__28522),
            .I(N__28519));
    LocalMux I__4720 (
            .O(N__28519),
            .I(N__28515));
    InMux I__4719 (
            .O(N__28518),
            .I(N__28512));
    Span4Mux_h I__4718 (
            .O(N__28515),
            .I(N__28506));
    LocalMux I__4717 (
            .O(N__28512),
            .I(N__28506));
    InMux I__4716 (
            .O(N__28511),
            .I(N__28503));
    Span4Mux_v I__4715 (
            .O(N__28506),
            .I(N__28500));
    LocalMux I__4714 (
            .O(N__28503),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__4713 (
            .O(N__28500),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__4712 (
            .O(N__28495),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__4711 (
            .O(N__28492),
            .I(N__28489));
    LocalMux I__4710 (
            .O(N__28489),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__4709 (
            .O(N__28486),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__4708 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__4707 (
            .O(N__28480),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__4706 (
            .O(N__28477),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__4705 (
            .O(N__28474),
            .I(N__28471));
    LocalMux I__4704 (
            .O(N__28471),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__4703 (
            .O(N__28468),
            .I(bfn_11_25_0_));
    InMux I__4702 (
            .O(N__28465),
            .I(N__28462));
    LocalMux I__4701 (
            .O(N__28462),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__4700 (
            .O(N__28459),
            .I(N__28456));
    LocalMux I__4699 (
            .O(N__28456),
            .I(N__28452));
    CascadeMux I__4698 (
            .O(N__28455),
            .I(N__28449));
    Span4Mux_h I__4697 (
            .O(N__28452),
            .I(N__28446));
    InMux I__4696 (
            .O(N__28449),
            .I(N__28442));
    Span4Mux_v I__4695 (
            .O(N__28446),
            .I(N__28439));
    InMux I__4694 (
            .O(N__28445),
            .I(N__28436));
    LocalMux I__4693 (
            .O(N__28442),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__4692 (
            .O(N__28439),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__4691 (
            .O(N__28436),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__4690 (
            .O(N__28429),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__4689 (
            .O(N__28426),
            .I(N__28423));
    LocalMux I__4688 (
            .O(N__28423),
            .I(N__28420));
    Span4Mux_v I__4687 (
            .O(N__28420),
            .I(N__28417));
    Odrv4 I__4686 (
            .O(N__28417),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__4685 (
            .O(N__28414),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__4684 (
            .O(N__28411),
            .I(N__28408));
    LocalMux I__4683 (
            .O(N__28408),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__4682 (
            .O(N__28405),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__4681 (
            .O(N__28402),
            .I(N__28399));
    LocalMux I__4680 (
            .O(N__28399),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__4679 (
            .O(N__28396),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__4678 (
            .O(N__28393),
            .I(N__28390));
    LocalMux I__4677 (
            .O(N__28390),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    CascadeMux I__4676 (
            .O(N__28387),
            .I(N__28384));
    InMux I__4675 (
            .O(N__28384),
            .I(N__28377));
    InMux I__4674 (
            .O(N__28383),
            .I(N__28377));
    CascadeMux I__4673 (
            .O(N__28382),
            .I(N__28374));
    LocalMux I__4672 (
            .O(N__28377),
            .I(N__28371));
    InMux I__4671 (
            .O(N__28374),
            .I(N__28368));
    Span4Mux_v I__4670 (
            .O(N__28371),
            .I(N__28365));
    LocalMux I__4669 (
            .O(N__28368),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__4668 (
            .O(N__28365),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__4667 (
            .O(N__28360),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__4666 (
            .O(N__28357),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__4665 (
            .O(N__28354),
            .I(N__28351));
    LocalMux I__4664 (
            .O(N__28351),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__4663 (
            .O(N__28348),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__4662 (
            .O(N__28345),
            .I(N__28342));
    LocalMux I__4661 (
            .O(N__28342),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__4660 (
            .O(N__28339),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__4659 (
            .O(N__28336),
            .I(N__28333));
    LocalMux I__4658 (
            .O(N__28333),
            .I(N__28330));
    Odrv12 I__4657 (
            .O(N__28330),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__4656 (
            .O(N__28327),
            .I(bfn_11_24_0_));
    InMux I__4655 (
            .O(N__28324),
            .I(N__28321));
    LocalMux I__4654 (
            .O(N__28321),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__4653 (
            .O(N__28318),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__4652 (
            .O(N__28315),
            .I(N__28312));
    LocalMux I__4651 (
            .O(N__28312),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__4650 (
            .O(N__28309),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__4649 (
            .O(N__28306),
            .I(N__28303));
    LocalMux I__4648 (
            .O(N__28303),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__4647 (
            .O(N__28300),
            .I(N__28296));
    InMux I__4646 (
            .O(N__28299),
            .I(N__28293));
    LocalMux I__4645 (
            .O(N__28296),
            .I(N__28290));
    LocalMux I__4644 (
            .O(N__28293),
            .I(N__28285));
    Span4Mux_v I__4643 (
            .O(N__28290),
            .I(N__28285));
    Span4Mux_v I__4642 (
            .O(N__28285),
            .I(N__28281));
    InMux I__4641 (
            .O(N__28284),
            .I(N__28278));
    Odrv4 I__4640 (
            .O(N__28281),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__4639 (
            .O(N__28278),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__4638 (
            .O(N__28273),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__4637 (
            .O(N__28270),
            .I(N__28267));
    LocalMux I__4636 (
            .O(N__28267),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__4635 (
            .O(N__28264),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__4634 (
            .O(N__28261),
            .I(N__28258));
    LocalMux I__4633 (
            .O(N__28258),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    CascadeMux I__4632 (
            .O(N__28255),
            .I(N__28251));
    CascadeMux I__4631 (
            .O(N__28254),
            .I(N__28248));
    InMux I__4630 (
            .O(N__28251),
            .I(N__28245));
    InMux I__4629 (
            .O(N__28248),
            .I(N__28242));
    LocalMux I__4628 (
            .O(N__28245),
            .I(N__28238));
    LocalMux I__4627 (
            .O(N__28242),
            .I(N__28235));
    InMux I__4626 (
            .O(N__28241),
            .I(N__28232));
    Span4Mux_h I__4625 (
            .O(N__28238),
            .I(N__28227));
    Span4Mux_v I__4624 (
            .O(N__28235),
            .I(N__28227));
    LocalMux I__4623 (
            .O(N__28232),
            .I(N__28224));
    Odrv4 I__4622 (
            .O(N__28227),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv12 I__4621 (
            .O(N__28224),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__4620 (
            .O(N__28219),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__4619 (
            .O(N__28216),
            .I(N__28213));
    LocalMux I__4618 (
            .O(N__28213),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__4617 (
            .O(N__28210),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__4616 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__4615 (
            .O(N__28204),
            .I(N__28201));
    Odrv4 I__4614 (
            .O(N__28201),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__4613 (
            .O(N__28198),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__4612 (
            .O(N__28195),
            .I(N__28192));
    LocalMux I__4611 (
            .O(N__28192),
            .I(N__28189));
    Odrv4 I__4610 (
            .O(N__28189),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__4609 (
            .O(N__28186),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__4608 (
            .O(N__28183),
            .I(N__28180));
    LocalMux I__4607 (
            .O(N__28180),
            .I(N__28177));
    Odrv4 I__4606 (
            .O(N__28177),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__4605 (
            .O(N__28174),
            .I(bfn_11_23_0_));
    InMux I__4604 (
            .O(N__28171),
            .I(N__28168));
    LocalMux I__4603 (
            .O(N__28168),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__4602 (
            .O(N__28165),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__4601 (
            .O(N__28162),
            .I(N__28159));
    LocalMux I__4600 (
            .O(N__28159),
            .I(N__28156));
    Span4Mux_h I__4599 (
            .O(N__28156),
            .I(N__28153));
    Odrv4 I__4598 (
            .O(N__28153),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__4597 (
            .O(N__28150),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__4596 (
            .O(N__28147),
            .I(N__28144));
    LocalMux I__4595 (
            .O(N__28144),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__4594 (
            .O(N__28141),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__4593 (
            .O(N__28138),
            .I(N__28135));
    LocalMux I__4592 (
            .O(N__28135),
            .I(N__28132));
    Span4Mux_h I__4591 (
            .O(N__28132),
            .I(N__28129));
    Odrv4 I__4590 (
            .O(N__28129),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__4589 (
            .O(N__28126),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__4588 (
            .O(N__28123),
            .I(N__28120));
    LocalMux I__4587 (
            .O(N__28120),
            .I(N__28117));
    Span4Mux_h I__4586 (
            .O(N__28117),
            .I(N__28114));
    Odrv4 I__4585 (
            .O(N__28114),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__4584 (
            .O(N__28111),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__4583 (
            .O(N__28108),
            .I(N__28105));
    LocalMux I__4582 (
            .O(N__28105),
            .I(N__28102));
    Span4Mux_h I__4581 (
            .O(N__28102),
            .I(N__28099));
    Span4Mux_v I__4580 (
            .O(N__28099),
            .I(N__28096));
    Odrv4 I__4579 (
            .O(N__28096),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__4578 (
            .O(N__28093),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__4577 (
            .O(N__28090),
            .I(N__28087));
    LocalMux I__4576 (
            .O(N__28087),
            .I(N__28084));
    Span4Mux_h I__4575 (
            .O(N__28084),
            .I(N__28081));
    Span4Mux_v I__4574 (
            .O(N__28081),
            .I(N__28078));
    Odrv4 I__4573 (
            .O(N__28078),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__4572 (
            .O(N__28075),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__4571 (
            .O(N__28072),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__4570 (
            .O(N__28069),
            .I(N__28066));
    LocalMux I__4569 (
            .O(N__28066),
            .I(N__28063));
    Span4Mux_v I__4568 (
            .O(N__28063),
            .I(N__28060));
    Odrv4 I__4567 (
            .O(N__28060),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__4566 (
            .O(N__28057),
            .I(N__28054));
    LocalMux I__4565 (
            .O(N__28054),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__4564 (
            .O(N__28051),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__4563 (
            .O(N__28048),
            .I(N__28045));
    LocalMux I__4562 (
            .O(N__28045),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__4561 (
            .O(N__28042),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__4560 (
            .O(N__28039),
            .I(N__28036));
    LocalMux I__4559 (
            .O(N__28036),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__4558 (
            .O(N__28033),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__4557 (
            .O(N__28030),
            .I(N__28027));
    LocalMux I__4556 (
            .O(N__28027),
            .I(N__28024));
    Span4Mux_h I__4555 (
            .O(N__28024),
            .I(N__28021));
    Sp12to4 I__4554 (
            .O(N__28021),
            .I(N__28018));
    Odrv12 I__4553 (
            .O(N__28018),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__4552 (
            .O(N__28015),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    CascadeMux I__4551 (
            .O(N__28012),
            .I(N__28009));
    InMux I__4550 (
            .O(N__28009),
            .I(N__28006));
    LocalMux I__4549 (
            .O(N__28006),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__4548 (
            .O(N__28003),
            .I(N__28000));
    LocalMux I__4547 (
            .O(N__28000),
            .I(N__27997));
    Span4Mux_h I__4546 (
            .O(N__27997),
            .I(N__27994));
    Odrv4 I__4545 (
            .O(N__27994),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__4544 (
            .O(N__27991),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__4543 (
            .O(N__27988),
            .I(N__27985));
    LocalMux I__4542 (
            .O(N__27985),
            .I(N__27982));
    Span4Mux_h I__4541 (
            .O(N__27982),
            .I(N__27979));
    Odrv4 I__4540 (
            .O(N__27979),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__4539 (
            .O(N__27976),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__4538 (
            .O(N__27973),
            .I(N__27970));
    InMux I__4537 (
            .O(N__27970),
            .I(N__27967));
    LocalMux I__4536 (
            .O(N__27967),
            .I(N__27964));
    Span12Mux_v I__4535 (
            .O(N__27964),
            .I(N__27961));
    Odrv12 I__4534 (
            .O(N__27961),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__4533 (
            .O(N__27958),
            .I(N__27955));
    LocalMux I__4532 (
            .O(N__27955),
            .I(N__27952));
    Span4Mux_v I__4531 (
            .O(N__27952),
            .I(N__27949));
    Odrv4 I__4530 (
            .O(N__27949),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__4529 (
            .O(N__27946),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__4528 (
            .O(N__27943),
            .I(N__27940));
    LocalMux I__4527 (
            .O(N__27940),
            .I(N__27937));
    Span12Mux_s11_h I__4526 (
            .O(N__27937),
            .I(N__27934));
    Odrv12 I__4525 (
            .O(N__27934),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__4524 (
            .O(N__27931),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__4523 (
            .O(N__27928),
            .I(N__27925));
    LocalMux I__4522 (
            .O(N__27925),
            .I(N__27922));
    Span4Mux_h I__4521 (
            .O(N__27922),
            .I(N__27919));
    Odrv4 I__4520 (
            .O(N__27919),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__4519 (
            .O(N__27916),
            .I(bfn_11_21_0_));
    InMux I__4518 (
            .O(N__27913),
            .I(N__27910));
    LocalMux I__4517 (
            .O(N__27910),
            .I(N__27907));
    Span4Mux_h I__4516 (
            .O(N__27907),
            .I(N__27904));
    Odrv4 I__4515 (
            .O(N__27904),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__4514 (
            .O(N__27901),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__4513 (
            .O(N__27898),
            .I(N__27895));
    InMux I__4512 (
            .O(N__27895),
            .I(N__27892));
    LocalMux I__4511 (
            .O(N__27892),
            .I(N__27889));
    Span4Mux_h I__4510 (
            .O(N__27889),
            .I(N__27886));
    Odrv4 I__4509 (
            .O(N__27886),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__4508 (
            .O(N__27883),
            .I(N__27880));
    LocalMux I__4507 (
            .O(N__27880),
            .I(N__27877));
    Span4Mux_h I__4506 (
            .O(N__27877),
            .I(N__27874));
    Odrv4 I__4505 (
            .O(N__27874),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__4504 (
            .O(N__27871),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__4503 (
            .O(N__27868),
            .I(N__27865));
    LocalMux I__4502 (
            .O(N__27865),
            .I(N__27862));
    Span4Mux_v I__4501 (
            .O(N__27862),
            .I(N__27859));
    Span4Mux_v I__4500 (
            .O(N__27859),
            .I(N__27856));
    Odrv4 I__4499 (
            .O(N__27856),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__4498 (
            .O(N__27853),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__4497 (
            .O(N__27850),
            .I(N__27847));
    LocalMux I__4496 (
            .O(N__27847),
            .I(N__27844));
    Span4Mux_h I__4495 (
            .O(N__27844),
            .I(N__27841));
    Sp12to4 I__4494 (
            .O(N__27841),
            .I(N__27838));
    Odrv12 I__4493 (
            .O(N__27838),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__4492 (
            .O(N__27835),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__4491 (
            .O(N__27832),
            .I(N__27829));
    LocalMux I__4490 (
            .O(N__27829),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__4489 (
            .O(N__27826),
            .I(N__27823));
    LocalMux I__4488 (
            .O(N__27823),
            .I(N__27820));
    Span4Mux_h I__4487 (
            .O(N__27820),
            .I(N__27817));
    Odrv4 I__4486 (
            .O(N__27817),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__4485 (
            .O(N__27814),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__4484 (
            .O(N__27811),
            .I(N__27808));
    LocalMux I__4483 (
            .O(N__27808),
            .I(N__27805));
    Span12Mux_v I__4482 (
            .O(N__27805),
            .I(N__27802));
    Odrv12 I__4481 (
            .O(N__27802),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__4480 (
            .O(N__27799),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__4479 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__4478 (
            .O(N__27793),
            .I(N__27790));
    Span4Mux_h I__4477 (
            .O(N__27790),
            .I(N__27787));
    Span4Mux_v I__4476 (
            .O(N__27787),
            .I(N__27784));
    Odrv4 I__4475 (
            .O(N__27784),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__4474 (
            .O(N__27781),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__4473 (
            .O(N__27778),
            .I(N__27775));
    LocalMux I__4472 (
            .O(N__27775),
            .I(N__27772));
    Span4Mux_v I__4471 (
            .O(N__27772),
            .I(N__27769));
    Span4Mux_v I__4470 (
            .O(N__27769),
            .I(N__27766));
    Odrv4 I__4469 (
            .O(N__27766),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__4468 (
            .O(N__27763),
            .I(bfn_11_20_0_));
    InMux I__4467 (
            .O(N__27760),
            .I(N__27757));
    LocalMux I__4466 (
            .O(N__27757),
            .I(N__27754));
    Span4Mux_v I__4465 (
            .O(N__27754),
            .I(N__27751));
    Span4Mux_v I__4464 (
            .O(N__27751),
            .I(N__27748));
    Span4Mux_h I__4463 (
            .O(N__27748),
            .I(N__27745));
    Odrv4 I__4462 (
            .O(N__27745),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__4461 (
            .O(N__27742),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__4460 (
            .O(N__27739),
            .I(N__27736));
    LocalMux I__4459 (
            .O(N__27736),
            .I(N__27733));
    Span4Mux_h I__4458 (
            .O(N__27733),
            .I(N__27730));
    Span4Mux_v I__4457 (
            .O(N__27730),
            .I(N__27727));
    Odrv4 I__4456 (
            .O(N__27727),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__4455 (
            .O(N__27724),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__4454 (
            .O(N__27721),
            .I(N__27718));
    LocalMux I__4453 (
            .O(N__27718),
            .I(N__27715));
    Span4Mux_h I__4452 (
            .O(N__27715),
            .I(N__27712));
    Span4Mux_v I__4451 (
            .O(N__27712),
            .I(N__27709));
    Odrv4 I__4450 (
            .O(N__27709),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__4449 (
            .O(N__27706),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__4448 (
            .O(N__27703),
            .I(N__27700));
    LocalMux I__4447 (
            .O(N__27700),
            .I(N__27697));
    Span4Mux_h I__4446 (
            .O(N__27697),
            .I(N__27694));
    Odrv4 I__4445 (
            .O(N__27694),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__4444 (
            .O(N__27691),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__4443 (
            .O(N__27688),
            .I(N__27685));
    LocalMux I__4442 (
            .O(N__27685),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__4441 (
            .O(N__27682),
            .I(N__27679));
    LocalMux I__4440 (
            .O(N__27679),
            .I(N__27676));
    Span4Mux_h I__4439 (
            .O(N__27676),
            .I(N__27673));
    Odrv4 I__4438 (
            .O(N__27673),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__4437 (
            .O(N__27670),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    InMux I__4436 (
            .O(N__27667),
            .I(N__27664));
    LocalMux I__4435 (
            .O(N__27664),
            .I(N__27661));
    Span12Mux_v I__4434 (
            .O(N__27661),
            .I(N__27658));
    Odrv12 I__4433 (
            .O(N__27658),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__4432 (
            .O(N__27655),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__4431 (
            .O(N__27652),
            .I(N__27649));
    LocalMux I__4430 (
            .O(N__27649),
            .I(N__27646));
    Span4Mux_h I__4429 (
            .O(N__27646),
            .I(N__27643));
    Span4Mux_v I__4428 (
            .O(N__27643),
            .I(N__27640));
    Odrv4 I__4427 (
            .O(N__27640),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__4426 (
            .O(N__27637),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__4425 (
            .O(N__27634),
            .I(N__27631));
    LocalMux I__4424 (
            .O(N__27631),
            .I(N__27628));
    Span4Mux_v I__4423 (
            .O(N__27628),
            .I(N__27625));
    Span4Mux_v I__4422 (
            .O(N__27625),
            .I(N__27622));
    Odrv4 I__4421 (
            .O(N__27622),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__4420 (
            .O(N__27619),
            .I(bfn_11_19_0_));
    InMux I__4419 (
            .O(N__27616),
            .I(N__27613));
    LocalMux I__4418 (
            .O(N__27613),
            .I(N__27610));
    Span4Mux_h I__4417 (
            .O(N__27610),
            .I(N__27607));
    Sp12to4 I__4416 (
            .O(N__27607),
            .I(N__27604));
    Span12Mux_v I__4415 (
            .O(N__27604),
            .I(N__27601));
    Odrv12 I__4414 (
            .O(N__27601),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__4413 (
            .O(N__27598),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__4412 (
            .O(N__27595),
            .I(N__27592));
    LocalMux I__4411 (
            .O(N__27592),
            .I(N__27589));
    Odrv4 I__4410 (
            .O(N__27589),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__4409 (
            .O(N__27586),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__4408 (
            .O(N__27583),
            .I(N__27580));
    LocalMux I__4407 (
            .O(N__27580),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__4406 (
            .O(N__27577),
            .I(N__27574));
    LocalMux I__4405 (
            .O(N__27574),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__4404 (
            .O(N__27571),
            .I(N__27568));
    LocalMux I__4403 (
            .O(N__27568),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__4402 (
            .O(N__27565),
            .I(N__27562));
    InMux I__4401 (
            .O(N__27562),
            .I(N__27559));
    LocalMux I__4400 (
            .O(N__27559),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__4399 (
            .O(N__27556),
            .I(N__27553));
    LocalMux I__4398 (
            .O(N__27553),
            .I(N__27550));
    Odrv4 I__4397 (
            .O(N__27550),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__4396 (
            .O(N__27547),
            .I(N__27544));
    InMux I__4395 (
            .O(N__27544),
            .I(N__27541));
    LocalMux I__4394 (
            .O(N__27541),
            .I(N__27538));
    Odrv4 I__4393 (
            .O(N__27538),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    CascadeMux I__4392 (
            .O(N__27535),
            .I(N__27532));
    InMux I__4391 (
            .O(N__27532),
            .I(N__27529));
    LocalMux I__4390 (
            .O(N__27529),
            .I(N__27526));
    Span4Mux_h I__4389 (
            .O(N__27526),
            .I(N__27522));
    InMux I__4388 (
            .O(N__27525),
            .I(N__27519));
    Span4Mux_v I__4387 (
            .O(N__27522),
            .I(N__27514));
    LocalMux I__4386 (
            .O(N__27519),
            .I(N__27514));
    Span4Mux_h I__4385 (
            .O(N__27514),
            .I(N__27511));
    Odrv4 I__4384 (
            .O(N__27511),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__4383 (
            .O(N__27508),
            .I(N__27505));
    InMux I__4382 (
            .O(N__27505),
            .I(N__27502));
    LocalMux I__4381 (
            .O(N__27502),
            .I(N__27498));
    InMux I__4380 (
            .O(N__27501),
            .I(N__27495));
    Span4Mux_v I__4379 (
            .O(N__27498),
            .I(N__27492));
    LocalMux I__4378 (
            .O(N__27495),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__4377 (
            .O(N__27492),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__4376 (
            .O(N__27487),
            .I(N__27484));
    InMux I__4375 (
            .O(N__27484),
            .I(N__27481));
    LocalMux I__4374 (
            .O(N__27481),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__4373 (
            .O(N__27478),
            .I(N__27475));
    LocalMux I__4372 (
            .O(N__27475),
            .I(N__27470));
    InMux I__4371 (
            .O(N__27474),
            .I(N__27466));
    InMux I__4370 (
            .O(N__27473),
            .I(N__27463));
    Span4Mux_h I__4369 (
            .O(N__27470),
            .I(N__27460));
    InMux I__4368 (
            .O(N__27469),
            .I(N__27457));
    LocalMux I__4367 (
            .O(N__27466),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__4366 (
            .O(N__27463),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__4365 (
            .O(N__27460),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__4364 (
            .O(N__27457),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    CascadeMux I__4363 (
            .O(N__27448),
            .I(N__27445));
    InMux I__4362 (
            .O(N__27445),
            .I(N__27442));
    LocalMux I__4361 (
            .O(N__27442),
            .I(N__27439));
    Odrv4 I__4360 (
            .O(N__27439),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__4359 (
            .O(N__27436),
            .I(N__27433));
    InMux I__4358 (
            .O(N__27433),
            .I(N__27430));
    LocalMux I__4357 (
            .O(N__27430),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    CascadeMux I__4356 (
            .O(N__27427),
            .I(N__27424));
    InMux I__4355 (
            .O(N__27424),
            .I(N__27421));
    LocalMux I__4354 (
            .O(N__27421),
            .I(N__27418));
    Odrv4 I__4353 (
            .O(N__27418),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__4352 (
            .O(N__27415),
            .I(N__27412));
    InMux I__4351 (
            .O(N__27412),
            .I(N__27408));
    InMux I__4350 (
            .O(N__27411),
            .I(N__27404));
    LocalMux I__4349 (
            .O(N__27408),
            .I(N__27401));
    CascadeMux I__4348 (
            .O(N__27407),
            .I(N__27398));
    LocalMux I__4347 (
            .O(N__27404),
            .I(N__27395));
    Span4Mux_h I__4346 (
            .O(N__27401),
            .I(N__27392));
    InMux I__4345 (
            .O(N__27398),
            .I(N__27389));
    Span4Mux_v I__4344 (
            .O(N__27395),
            .I(N__27386));
    Span4Mux_v I__4343 (
            .O(N__27392),
            .I(N__27382));
    LocalMux I__4342 (
            .O(N__27389),
            .I(N__27377));
    Span4Mux_h I__4341 (
            .O(N__27386),
            .I(N__27377));
    InMux I__4340 (
            .O(N__27385),
            .I(N__27374));
    Odrv4 I__4339 (
            .O(N__27382),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__4338 (
            .O(N__27377),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__4337 (
            .O(N__27374),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__4336 (
            .O(N__27367),
            .I(N__27364));
    InMux I__4335 (
            .O(N__27364),
            .I(N__27361));
    LocalMux I__4334 (
            .O(N__27361),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__4333 (
            .O(N__27358),
            .I(N__27355));
    InMux I__4332 (
            .O(N__27355),
            .I(N__27352));
    LocalMux I__4331 (
            .O(N__27352),
            .I(N__27349));
    Odrv4 I__4330 (
            .O(N__27349),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__4329 (
            .O(N__27346),
            .I(N__27343));
    LocalMux I__4328 (
            .O(N__27343),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__4327 (
            .O(N__27340),
            .I(N__27337));
    LocalMux I__4326 (
            .O(N__27337),
            .I(N__27334));
    Span4Mux_h I__4325 (
            .O(N__27334),
            .I(N__27331));
    Span4Mux_v I__4324 (
            .O(N__27331),
            .I(N__27326));
    InMux I__4323 (
            .O(N__27330),
            .I(N__27323));
    InMux I__4322 (
            .O(N__27329),
            .I(N__27319));
    Span4Mux_h I__4321 (
            .O(N__27326),
            .I(N__27314));
    LocalMux I__4320 (
            .O(N__27323),
            .I(N__27314));
    InMux I__4319 (
            .O(N__27322),
            .I(N__27311));
    LocalMux I__4318 (
            .O(N__27319),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__4317 (
            .O(N__27314),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__4316 (
            .O(N__27311),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__4315 (
            .O(N__27304),
            .I(N__27301));
    InMux I__4314 (
            .O(N__27301),
            .I(N__27298));
    LocalMux I__4313 (
            .O(N__27298),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__4312 (
            .O(N__27295),
            .I(N__27292));
    InMux I__4311 (
            .O(N__27292),
            .I(N__27289));
    LocalMux I__4310 (
            .O(N__27289),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__4309 (
            .O(N__27286),
            .I(N__27283));
    LocalMux I__4308 (
            .O(N__27283),
            .I(N__27278));
    InMux I__4307 (
            .O(N__27282),
            .I(N__27273));
    InMux I__4306 (
            .O(N__27281),
            .I(N__27273));
    Span4Mux_v I__4305 (
            .O(N__27278),
            .I(N__27268));
    LocalMux I__4304 (
            .O(N__27273),
            .I(N__27268));
    Span4Mux_h I__4303 (
            .O(N__27268),
            .I(N__27264));
    InMux I__4302 (
            .O(N__27267),
            .I(N__27261));
    Odrv4 I__4301 (
            .O(N__27264),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__4300 (
            .O(N__27261),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__4299 (
            .O(N__27256),
            .I(N__27253));
    LocalMux I__4298 (
            .O(N__27253),
            .I(N__27249));
    InMux I__4297 (
            .O(N__27252),
            .I(N__27246));
    Odrv4 I__4296 (
            .O(N__27249),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__4295 (
            .O(N__27246),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__4294 (
            .O(N__27241),
            .I(N__27235));
    InMux I__4293 (
            .O(N__27240),
            .I(N__27235));
    LocalMux I__4292 (
            .O(N__27235),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__4291 (
            .O(N__27232),
            .I(N__27227));
    InMux I__4290 (
            .O(N__27231),
            .I(N__27224));
    InMux I__4289 (
            .O(N__27230),
            .I(N__27221));
    LocalMux I__4288 (
            .O(N__27227),
            .I(N__27218));
    LocalMux I__4287 (
            .O(N__27224),
            .I(N__27215));
    LocalMux I__4286 (
            .O(N__27221),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv12 I__4285 (
            .O(N__27218),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv4 I__4284 (
            .O(N__27215),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__4283 (
            .O(N__27208),
            .I(N__27203));
    InMux I__4282 (
            .O(N__27207),
            .I(N__27200));
    InMux I__4281 (
            .O(N__27206),
            .I(N__27197));
    LocalMux I__4280 (
            .O(N__27203),
            .I(N__27194));
    LocalMux I__4279 (
            .O(N__27200),
            .I(N__27191));
    LocalMux I__4278 (
            .O(N__27197),
            .I(N__27188));
    Span4Mux_v I__4277 (
            .O(N__27194),
            .I(N__27184));
    Span4Mux_h I__4276 (
            .O(N__27191),
            .I(N__27179));
    Span4Mux_h I__4275 (
            .O(N__27188),
            .I(N__27179));
    InMux I__4274 (
            .O(N__27187),
            .I(N__27176));
    Odrv4 I__4273 (
            .O(N__27184),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__4272 (
            .O(N__27179),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__4271 (
            .O(N__27176),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    CascadeMux I__4270 (
            .O(N__27169),
            .I(N__27166));
    InMux I__4269 (
            .O(N__27166),
            .I(N__27160));
    InMux I__4268 (
            .O(N__27165),
            .I(N__27160));
    LocalMux I__4267 (
            .O(N__27160),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__4266 (
            .O(N__27157),
            .I(N__27154));
    InMux I__4265 (
            .O(N__27154),
            .I(N__27148));
    InMux I__4264 (
            .O(N__27153),
            .I(N__27145));
    InMux I__4263 (
            .O(N__27152),
            .I(N__27140));
    InMux I__4262 (
            .O(N__27151),
            .I(N__27140));
    LocalMux I__4261 (
            .O(N__27148),
            .I(N__27135));
    LocalMux I__4260 (
            .O(N__27145),
            .I(N__27135));
    LocalMux I__4259 (
            .O(N__27140),
            .I(N__27132));
    Span4Mux_v I__4258 (
            .O(N__27135),
            .I(N__27129));
    Span4Mux_h I__4257 (
            .O(N__27132),
            .I(N__27126));
    Odrv4 I__4256 (
            .O(N__27129),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__4255 (
            .O(N__27126),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__4254 (
            .O(N__27121),
            .I(N__27118));
    LocalMux I__4253 (
            .O(N__27118),
            .I(N__27113));
    InMux I__4252 (
            .O(N__27117),
            .I(N__27110));
    InMux I__4251 (
            .O(N__27116),
            .I(N__27107));
    Span4Mux_v I__4250 (
            .O(N__27113),
            .I(N__27104));
    LocalMux I__4249 (
            .O(N__27110),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__4248 (
            .O(N__27107),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__4247 (
            .O(N__27104),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    InMux I__4246 (
            .O(N__27097),
            .I(N__27091));
    InMux I__4245 (
            .O(N__27096),
            .I(N__27091));
    LocalMux I__4244 (
            .O(N__27091),
            .I(N__27088));
    Odrv12 I__4243 (
            .O(N__27088),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    InMux I__4242 (
            .O(N__27085),
            .I(N__27082));
    LocalMux I__4241 (
            .O(N__27082),
            .I(N__27077));
    InMux I__4240 (
            .O(N__27081),
            .I(N__27074));
    InMux I__4239 (
            .O(N__27080),
            .I(N__27071));
    Span4Mux_h I__4238 (
            .O(N__27077),
            .I(N__27068));
    LocalMux I__4237 (
            .O(N__27074),
            .I(N__27065));
    LocalMux I__4236 (
            .O(N__27071),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__4235 (
            .O(N__27068),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv12 I__4234 (
            .O(N__27065),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__4233 (
            .O(N__27058),
            .I(N__27054));
    InMux I__4232 (
            .O(N__27057),
            .I(N__27050));
    LocalMux I__4231 (
            .O(N__27054),
            .I(N__27047));
    InMux I__4230 (
            .O(N__27053),
            .I(N__27044));
    LocalMux I__4229 (
            .O(N__27050),
            .I(N__27041));
    Span4Mux_v I__4228 (
            .O(N__27047),
            .I(N__27037));
    LocalMux I__4227 (
            .O(N__27044),
            .I(N__27034));
    Span4Mux_v I__4226 (
            .O(N__27041),
            .I(N__27031));
    InMux I__4225 (
            .O(N__27040),
            .I(N__27028));
    Odrv4 I__4224 (
            .O(N__27037),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__4223 (
            .O(N__27034),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__4222 (
            .O(N__27031),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__4221 (
            .O(N__27028),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__4220 (
            .O(N__27019),
            .I(N__27016));
    InMux I__4219 (
            .O(N__27016),
            .I(N__27010));
    InMux I__4218 (
            .O(N__27015),
            .I(N__27010));
    LocalMux I__4217 (
            .O(N__27010),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    InMux I__4216 (
            .O(N__27007),
            .I(N__27003));
    InMux I__4215 (
            .O(N__27006),
            .I(N__26998));
    LocalMux I__4214 (
            .O(N__27003),
            .I(N__26995));
    InMux I__4213 (
            .O(N__27002),
            .I(N__26990));
    InMux I__4212 (
            .O(N__27001),
            .I(N__26990));
    LocalMux I__4211 (
            .O(N__26998),
            .I(N__26987));
    Span4Mux_h I__4210 (
            .O(N__26995),
            .I(N__26982));
    LocalMux I__4209 (
            .O(N__26990),
            .I(N__26982));
    Span4Mux_h I__4208 (
            .O(N__26987),
            .I(N__26979));
    Span4Mux_v I__4207 (
            .O(N__26982),
            .I(N__26976));
    Odrv4 I__4206 (
            .O(N__26979),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__4205 (
            .O(N__26976),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__4204 (
            .O(N__26971),
            .I(N__26968));
    LocalMux I__4203 (
            .O(N__26968),
            .I(N__26964));
    InMux I__4202 (
            .O(N__26967),
            .I(N__26960));
    Span12Mux_h I__4201 (
            .O(N__26964),
            .I(N__26957));
    InMux I__4200 (
            .O(N__26963),
            .I(N__26954));
    LocalMux I__4199 (
            .O(N__26960),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv12 I__4198 (
            .O(N__26957),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__4197 (
            .O(N__26954),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__4196 (
            .O(N__26947),
            .I(N__26944));
    LocalMux I__4195 (
            .O(N__26944),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__4194 (
            .O(N__26941),
            .I(N__26938));
    LocalMux I__4193 (
            .O(N__26938),
            .I(N__26935));
    Span4Mux_h I__4192 (
            .O(N__26935),
            .I(N__26931));
    InMux I__4191 (
            .O(N__26934),
            .I(N__26927));
    Span4Mux_v I__4190 (
            .O(N__26931),
            .I(N__26924));
    InMux I__4189 (
            .O(N__26930),
            .I(N__26921));
    LocalMux I__4188 (
            .O(N__26927),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__4187 (
            .O(N__26924),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__4186 (
            .O(N__26921),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__4185 (
            .O(N__26914),
            .I(N__26908));
    InMux I__4184 (
            .O(N__26913),
            .I(N__26905));
    InMux I__4183 (
            .O(N__26912),
            .I(N__26902));
    InMux I__4182 (
            .O(N__26911),
            .I(N__26899));
    LocalMux I__4181 (
            .O(N__26908),
            .I(N__26896));
    LocalMux I__4180 (
            .O(N__26905),
            .I(N__26893));
    LocalMux I__4179 (
            .O(N__26902),
            .I(N__26890));
    LocalMux I__4178 (
            .O(N__26899),
            .I(N__26887));
    Span4Mux_v I__4177 (
            .O(N__26896),
            .I(N__26880));
    Span4Mux_h I__4176 (
            .O(N__26893),
            .I(N__26880));
    Span4Mux_h I__4175 (
            .O(N__26890),
            .I(N__26880));
    Odrv12 I__4174 (
            .O(N__26887),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__4173 (
            .O(N__26880),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__4172 (
            .O(N__26875),
            .I(N__26869));
    InMux I__4171 (
            .O(N__26874),
            .I(N__26869));
    LocalMux I__4170 (
            .O(N__26869),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__4169 (
            .O(N__26866),
            .I(N__26862));
    CascadeMux I__4168 (
            .O(N__26865),
            .I(N__26857));
    LocalMux I__4167 (
            .O(N__26862),
            .I(N__26854));
    InMux I__4166 (
            .O(N__26861),
            .I(N__26849));
    InMux I__4165 (
            .O(N__26860),
            .I(N__26849));
    InMux I__4164 (
            .O(N__26857),
            .I(N__26846));
    Span4Mux_h I__4163 (
            .O(N__26854),
            .I(N__26843));
    LocalMux I__4162 (
            .O(N__26849),
            .I(N__26840));
    LocalMux I__4161 (
            .O(N__26846),
            .I(N__26837));
    Odrv4 I__4160 (
            .O(N__26843),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv12 I__4159 (
            .O(N__26840),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__4158 (
            .O(N__26837),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__4157 (
            .O(N__26830),
            .I(N__26827));
    LocalMux I__4156 (
            .O(N__26827),
            .I(N__26824));
    Span4Mux_v I__4155 (
            .O(N__26824),
            .I(N__26821));
    Span4Mux_h I__4154 (
            .O(N__26821),
            .I(N__26817));
    InMux I__4153 (
            .O(N__26820),
            .I(N__26814));
    Odrv4 I__4152 (
            .O(N__26817),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__4151 (
            .O(N__26814),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__4150 (
            .O(N__26809),
            .I(N__26806));
    InMux I__4149 (
            .O(N__26806),
            .I(N__26800));
    InMux I__4148 (
            .O(N__26805),
            .I(N__26800));
    LocalMux I__4147 (
            .O(N__26800),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__4146 (
            .O(N__26797),
            .I(N__26794));
    LocalMux I__4145 (
            .O(N__26794),
            .I(N__26788));
    InMux I__4144 (
            .O(N__26793),
            .I(N__26783));
    InMux I__4143 (
            .O(N__26792),
            .I(N__26783));
    InMux I__4142 (
            .O(N__26791),
            .I(N__26780));
    Span4Mux_h I__4141 (
            .O(N__26788),
            .I(N__26777));
    LocalMux I__4140 (
            .O(N__26783),
            .I(N__26774));
    LocalMux I__4139 (
            .O(N__26780),
            .I(N__26771));
    Odrv4 I__4138 (
            .O(N__26777),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__4137 (
            .O(N__26774),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__4136 (
            .O(N__26771),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__4135 (
            .O(N__26764),
            .I(N__26761));
    LocalMux I__4134 (
            .O(N__26761),
            .I(N__26758));
    Span4Mux_v I__4133 (
            .O(N__26758),
            .I(N__26755));
    Span4Mux_h I__4132 (
            .O(N__26755),
            .I(N__26751));
    InMux I__4131 (
            .O(N__26754),
            .I(N__26748));
    Odrv4 I__4130 (
            .O(N__26751),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__4129 (
            .O(N__26748),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__4128 (
            .O(N__26743),
            .I(N__26737));
    InMux I__4127 (
            .O(N__26742),
            .I(N__26737));
    LocalMux I__4126 (
            .O(N__26737),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__4125 (
            .O(N__26734),
            .I(N__26731));
    LocalMux I__4124 (
            .O(N__26731),
            .I(N__26728));
    Span4Mux_h I__4123 (
            .O(N__26728),
            .I(N__26723));
    InMux I__4122 (
            .O(N__26727),
            .I(N__26720));
    InMux I__4121 (
            .O(N__26726),
            .I(N__26717));
    Span4Mux_v I__4120 (
            .O(N__26723),
            .I(N__26714));
    LocalMux I__4119 (
            .O(N__26720),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__4118 (
            .O(N__26717),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__4117 (
            .O(N__26714),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    InMux I__4116 (
            .O(N__26707),
            .I(N__26702));
    InMux I__4115 (
            .O(N__26706),
            .I(N__26699));
    InMux I__4114 (
            .O(N__26705),
            .I(N__26696));
    LocalMux I__4113 (
            .O(N__26702),
            .I(N__26693));
    LocalMux I__4112 (
            .O(N__26699),
            .I(N__26690));
    LocalMux I__4111 (
            .O(N__26696),
            .I(N__26687));
    Span4Mux_h I__4110 (
            .O(N__26693),
            .I(N__26683));
    Span4Mux_h I__4109 (
            .O(N__26690),
            .I(N__26678));
    Span4Mux_h I__4108 (
            .O(N__26687),
            .I(N__26678));
    InMux I__4107 (
            .O(N__26686),
            .I(N__26675));
    Odrv4 I__4106 (
            .O(N__26683),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__4105 (
            .O(N__26678),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__4104 (
            .O(N__26675),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__4103 (
            .O(N__26668),
            .I(N__26665));
    InMux I__4102 (
            .O(N__26665),
            .I(N__26659));
    InMux I__4101 (
            .O(N__26664),
            .I(N__26659));
    LocalMux I__4100 (
            .O(N__26659),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__4099 (
            .O(N__26656),
            .I(N__26653));
    LocalMux I__4098 (
            .O(N__26653),
            .I(N__26649));
    InMux I__4097 (
            .O(N__26652),
            .I(N__26646));
    Span4Mux_v I__4096 (
            .O(N__26649),
            .I(N__26640));
    LocalMux I__4095 (
            .O(N__26646),
            .I(N__26640));
    InMux I__4094 (
            .O(N__26645),
            .I(N__26637));
    Span4Mux_h I__4093 (
            .O(N__26640),
            .I(N__26634));
    LocalMux I__4092 (
            .O(N__26637),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__4091 (
            .O(N__26634),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__4090 (
            .O(N__26629),
            .I(N__26625));
    InMux I__4089 (
            .O(N__26628),
            .I(N__26622));
    LocalMux I__4088 (
            .O(N__26625),
            .I(N__26617));
    LocalMux I__4087 (
            .O(N__26622),
            .I(N__26617));
    Span4Mux_v I__4086 (
            .O(N__26617),
            .I(N__26612));
    InMux I__4085 (
            .O(N__26616),
            .I(N__26607));
    InMux I__4084 (
            .O(N__26615),
            .I(N__26607));
    Odrv4 I__4083 (
            .O(N__26612),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__4082 (
            .O(N__26607),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__4081 (
            .O(N__26602),
            .I(N__26598));
    InMux I__4080 (
            .O(N__26601),
            .I(N__26595));
    LocalMux I__4079 (
            .O(N__26598),
            .I(N__26590));
    LocalMux I__4078 (
            .O(N__26595),
            .I(N__26587));
    InMux I__4077 (
            .O(N__26594),
            .I(N__26584));
    InMux I__4076 (
            .O(N__26593),
            .I(N__26581));
    Span4Mux_h I__4075 (
            .O(N__26590),
            .I(N__26578));
    Span4Mux_h I__4074 (
            .O(N__26587),
            .I(N__26575));
    LocalMux I__4073 (
            .O(N__26584),
            .I(N__26570));
    LocalMux I__4072 (
            .O(N__26581),
            .I(N__26570));
    Odrv4 I__4071 (
            .O(N__26578),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__4070 (
            .O(N__26575),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__4069 (
            .O(N__26570),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__4068 (
            .O(N__26563),
            .I(N__26560));
    LocalMux I__4067 (
            .O(N__26560),
            .I(N__26556));
    InMux I__4066 (
            .O(N__26559),
            .I(N__26552));
    Span4Mux_v I__4065 (
            .O(N__26556),
            .I(N__26549));
    InMux I__4064 (
            .O(N__26555),
            .I(N__26546));
    LocalMux I__4063 (
            .O(N__26552),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__4062 (
            .O(N__26549),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__4061 (
            .O(N__26546),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__4060 (
            .O(N__26539),
            .I(N__26534));
    InMux I__4059 (
            .O(N__26538),
            .I(N__26531));
    InMux I__4058 (
            .O(N__26537),
            .I(N__26528));
    LocalMux I__4057 (
            .O(N__26534),
            .I(N__26525));
    LocalMux I__4056 (
            .O(N__26531),
            .I(N__26520));
    LocalMux I__4055 (
            .O(N__26528),
            .I(N__26520));
    Span4Mux_v I__4054 (
            .O(N__26525),
            .I(N__26514));
    Span4Mux_v I__4053 (
            .O(N__26520),
            .I(N__26514));
    InMux I__4052 (
            .O(N__26519),
            .I(N__26511));
    Odrv4 I__4051 (
            .O(N__26514),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__4050 (
            .O(N__26511),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__4049 (
            .O(N__26506),
            .I(N__26503));
    LocalMux I__4048 (
            .O(N__26503),
            .I(N__26499));
    InMux I__4047 (
            .O(N__26502),
            .I(N__26496));
    Odrv4 I__4046 (
            .O(N__26499),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    LocalMux I__4045 (
            .O(N__26496),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__4044 (
            .O(N__26491),
            .I(N__26486));
    InMux I__4043 (
            .O(N__26490),
            .I(N__26481));
    InMux I__4042 (
            .O(N__26489),
            .I(N__26481));
    LocalMux I__4041 (
            .O(N__26486),
            .I(N__26475));
    LocalMux I__4040 (
            .O(N__26481),
            .I(N__26475));
    CascadeMux I__4039 (
            .O(N__26480),
            .I(N__26472));
    Span4Mux_v I__4038 (
            .O(N__26475),
            .I(N__26469));
    InMux I__4037 (
            .O(N__26472),
            .I(N__26466));
    Odrv4 I__4036 (
            .O(N__26469),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__4035 (
            .O(N__26466),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__4034 (
            .O(N__26461),
            .I(N__26456));
    InMux I__4033 (
            .O(N__26460),
            .I(N__26453));
    InMux I__4032 (
            .O(N__26459),
            .I(N__26449));
    LocalMux I__4031 (
            .O(N__26456),
            .I(N__26446));
    LocalMux I__4030 (
            .O(N__26453),
            .I(N__26443));
    InMux I__4029 (
            .O(N__26452),
            .I(N__26440));
    LocalMux I__4028 (
            .O(N__26449),
            .I(N__26437));
    Span12Mux_h I__4027 (
            .O(N__26446),
            .I(N__26434));
    Span4Mux_h I__4026 (
            .O(N__26443),
            .I(N__26431));
    LocalMux I__4025 (
            .O(N__26440),
            .I(N__26428));
    Span4Mux_h I__4024 (
            .O(N__26437),
            .I(N__26425));
    Odrv12 I__4023 (
            .O(N__26434),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__4022 (
            .O(N__26431),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__4021 (
            .O(N__26428),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__4020 (
            .O(N__26425),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__4019 (
            .O(N__26416),
            .I(N__26413));
    LocalMux I__4018 (
            .O(N__26413),
            .I(N__26410));
    Span4Mux_h I__4017 (
            .O(N__26410),
            .I(N__26406));
    InMux I__4016 (
            .O(N__26409),
            .I(N__26402));
    Span4Mux_v I__4015 (
            .O(N__26406),
            .I(N__26399));
    InMux I__4014 (
            .O(N__26405),
            .I(N__26396));
    LocalMux I__4013 (
            .O(N__26402),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv4 I__4012 (
            .O(N__26399),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__4011 (
            .O(N__26396),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    CascadeMux I__4010 (
            .O(N__26389),
            .I(N__26384));
    InMux I__4009 (
            .O(N__26388),
            .I(N__26381));
    InMux I__4008 (
            .O(N__26387),
            .I(N__26375));
    InMux I__4007 (
            .O(N__26384),
            .I(N__26375));
    LocalMux I__4006 (
            .O(N__26381),
            .I(N__26372));
    InMux I__4005 (
            .O(N__26380),
            .I(N__26369));
    LocalMux I__4004 (
            .O(N__26375),
            .I(N__26366));
    Span4Mux_h I__4003 (
            .O(N__26372),
            .I(N__26363));
    LocalMux I__4002 (
            .O(N__26369),
            .I(N__26360));
    Span4Mux_h I__4001 (
            .O(N__26366),
            .I(N__26357));
    Odrv4 I__4000 (
            .O(N__26363),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__3999 (
            .O(N__26360),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__3998 (
            .O(N__26357),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__3997 (
            .O(N__26350),
            .I(N__26346));
    InMux I__3996 (
            .O(N__26349),
            .I(N__26343));
    LocalMux I__3995 (
            .O(N__26346),
            .I(N__26337));
    LocalMux I__3994 (
            .O(N__26343),
            .I(N__26337));
    InMux I__3993 (
            .O(N__26342),
            .I(N__26334));
    Span12Mux_s11_v I__3992 (
            .O(N__26337),
            .I(N__26331));
    LocalMux I__3991 (
            .O(N__26334),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv12 I__3990 (
            .O(N__26331),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__3989 (
            .O(N__26326),
            .I(N__26323));
    LocalMux I__3988 (
            .O(N__26323),
            .I(N__26317));
    InMux I__3987 (
            .O(N__26322),
            .I(N__26312));
    InMux I__3986 (
            .O(N__26321),
            .I(N__26312));
    InMux I__3985 (
            .O(N__26320),
            .I(N__26309));
    Odrv4 I__3984 (
            .O(N__26317),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__3983 (
            .O(N__26312),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__3982 (
            .O(N__26309),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__3981 (
            .O(N__26302),
            .I(N__26299));
    LocalMux I__3980 (
            .O(N__26299),
            .I(N__26295));
    InMux I__3979 (
            .O(N__26298),
            .I(N__26292));
    Odrv4 I__3978 (
            .O(N__26295),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__3977 (
            .O(N__26292),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__3976 (
            .O(N__26287),
            .I(N__26281));
    InMux I__3975 (
            .O(N__26286),
            .I(N__26276));
    InMux I__3974 (
            .O(N__26285),
            .I(N__26276));
    InMux I__3973 (
            .O(N__26284),
            .I(N__26273));
    LocalMux I__3972 (
            .O(N__26281),
            .I(N__26268));
    LocalMux I__3971 (
            .O(N__26276),
            .I(N__26268));
    LocalMux I__3970 (
            .O(N__26273),
            .I(N__26265));
    Span4Mux_v I__3969 (
            .O(N__26268),
            .I(N__26260));
    Span4Mux_v I__3968 (
            .O(N__26265),
            .I(N__26260));
    Odrv4 I__3967 (
            .O(N__26260),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__3966 (
            .O(N__26257),
            .I(N__26253));
    InMux I__3965 (
            .O(N__26256),
            .I(N__26250));
    LocalMux I__3964 (
            .O(N__26253),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__3963 (
            .O(N__26250),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    CascadeMux I__3962 (
            .O(N__26245),
            .I(N__26242));
    InMux I__3961 (
            .O(N__26242),
            .I(N__26239));
    LocalMux I__3960 (
            .O(N__26239),
            .I(N__26236));
    Odrv4 I__3959 (
            .O(N__26236),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__3958 (
            .O(N__26233),
            .I(N__26226));
    InMux I__3957 (
            .O(N__26232),
            .I(N__26226));
    InMux I__3956 (
            .O(N__26231),
            .I(N__26223));
    LocalMux I__3955 (
            .O(N__26226),
            .I(N__26220));
    LocalMux I__3954 (
            .O(N__26223),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__3953 (
            .O(N__26220),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__3952 (
            .O(N__26215),
            .I(N__26212));
    InMux I__3951 (
            .O(N__26212),
            .I(N__26205));
    InMux I__3950 (
            .O(N__26211),
            .I(N__26205));
    InMux I__3949 (
            .O(N__26210),
            .I(N__26202));
    LocalMux I__3948 (
            .O(N__26205),
            .I(N__26199));
    LocalMux I__3947 (
            .O(N__26202),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv12 I__3946 (
            .O(N__26199),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__3945 (
            .O(N__26194),
            .I(N__26191));
    LocalMux I__3944 (
            .O(N__26191),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    CascadeMux I__3943 (
            .O(N__26188),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__3942 (
            .O(N__26185),
            .I(N__26182));
    LocalMux I__3941 (
            .O(N__26182),
            .I(N__26179));
    Span4Mux_h I__3940 (
            .O(N__26179),
            .I(N__26176));
    Odrv4 I__3939 (
            .O(N__26176),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__3938 (
            .O(N__26173),
            .I(N__26170));
    LocalMux I__3937 (
            .O(N__26170),
            .I(N__26166));
    InMux I__3936 (
            .O(N__26169),
            .I(N__26163));
    Span4Mux_v I__3935 (
            .O(N__26166),
            .I(N__26159));
    LocalMux I__3934 (
            .O(N__26163),
            .I(N__26156));
    InMux I__3933 (
            .O(N__26162),
            .I(N__26153));
    Span4Mux_h I__3932 (
            .O(N__26159),
            .I(N__26148));
    Span4Mux_h I__3931 (
            .O(N__26156),
            .I(N__26148));
    LocalMux I__3930 (
            .O(N__26153),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv4 I__3929 (
            .O(N__26148),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    InMux I__3928 (
            .O(N__26143),
            .I(N__26138));
    InMux I__3927 (
            .O(N__26142),
            .I(N__26135));
    InMux I__3926 (
            .O(N__26141),
            .I(N__26132));
    LocalMux I__3925 (
            .O(N__26138),
            .I(N__26128));
    LocalMux I__3924 (
            .O(N__26135),
            .I(N__26125));
    LocalMux I__3923 (
            .O(N__26132),
            .I(N__26122));
    CascadeMux I__3922 (
            .O(N__26131),
            .I(N__26119));
    Span4Mux_v I__3921 (
            .O(N__26128),
            .I(N__26114));
    Span4Mux_v I__3920 (
            .O(N__26125),
            .I(N__26114));
    Span4Mux_h I__3919 (
            .O(N__26122),
            .I(N__26111));
    InMux I__3918 (
            .O(N__26119),
            .I(N__26108));
    Odrv4 I__3917 (
            .O(N__26114),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv4 I__3916 (
            .O(N__26111),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__3915 (
            .O(N__26108),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    CascadeMux I__3914 (
            .O(N__26101),
            .I(N__26098));
    InMux I__3913 (
            .O(N__26098),
            .I(N__26092));
    InMux I__3912 (
            .O(N__26097),
            .I(N__26092));
    LocalMux I__3911 (
            .O(N__26092),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    CascadeMux I__3910 (
            .O(N__26089),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__3909 (
            .O(N__26086),
            .I(N__26080));
    InMux I__3908 (
            .O(N__26085),
            .I(N__26080));
    LocalMux I__3907 (
            .O(N__26080),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__3906 (
            .O(N__26077),
            .I(N__26073));
    InMux I__3905 (
            .O(N__26076),
            .I(N__26069));
    LocalMux I__3904 (
            .O(N__26073),
            .I(N__26065));
    InMux I__3903 (
            .O(N__26072),
            .I(N__26062));
    LocalMux I__3902 (
            .O(N__26069),
            .I(N__26059));
    InMux I__3901 (
            .O(N__26068),
            .I(N__26056));
    Span4Mux_v I__3900 (
            .O(N__26065),
            .I(N__26053));
    LocalMux I__3899 (
            .O(N__26062),
            .I(N__26050));
    Span4Mux_h I__3898 (
            .O(N__26059),
            .I(N__26045));
    LocalMux I__3897 (
            .O(N__26056),
            .I(N__26045));
    Odrv4 I__3896 (
            .O(N__26053),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv12 I__3895 (
            .O(N__26050),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__3894 (
            .O(N__26045),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__3893 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__3892 (
            .O(N__26035),
            .I(N__26031));
    InMux I__3891 (
            .O(N__26034),
            .I(N__26027));
    Span4Mux_v I__3890 (
            .O(N__26031),
            .I(N__26024));
    InMux I__3889 (
            .O(N__26030),
            .I(N__26021));
    LocalMux I__3888 (
            .O(N__26027),
            .I(N__26018));
    Span4Mux_h I__3887 (
            .O(N__26024),
            .I(N__26015));
    LocalMux I__3886 (
            .O(N__26021),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv4 I__3885 (
            .O(N__26018),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv4 I__3884 (
            .O(N__26015),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__3883 (
            .O(N__26008),
            .I(N__26005));
    LocalMux I__3882 (
            .O(N__26005),
            .I(N__26002));
    Span4Mux_h I__3881 (
            .O(N__26002),
            .I(N__25998));
    InMux I__3880 (
            .O(N__26001),
            .I(N__25995));
    Span4Mux_v I__3879 (
            .O(N__25998),
            .I(N__25989));
    LocalMux I__3878 (
            .O(N__25995),
            .I(N__25989));
    InMux I__3877 (
            .O(N__25994),
            .I(N__25986));
    Span4Mux_h I__3876 (
            .O(N__25989),
            .I(N__25983));
    LocalMux I__3875 (
            .O(N__25986),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__3874 (
            .O(N__25983),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    CascadeMux I__3873 (
            .O(N__25978),
            .I(N__25975));
    InMux I__3872 (
            .O(N__25975),
            .I(N__25972));
    LocalMux I__3871 (
            .O(N__25972),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__3870 (
            .O(N__25969),
            .I(N__25966));
    LocalMux I__3869 (
            .O(N__25966),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__3868 (
            .O(N__25963),
            .I(N__25960));
    InMux I__3867 (
            .O(N__25960),
            .I(N__25957));
    LocalMux I__3866 (
            .O(N__25957),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__3865 (
            .O(N__25954),
            .I(N__25947));
    InMux I__3864 (
            .O(N__25953),
            .I(N__25947));
    InMux I__3863 (
            .O(N__25952),
            .I(N__25944));
    LocalMux I__3862 (
            .O(N__25947),
            .I(N__25941));
    LocalMux I__3861 (
            .O(N__25944),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__3860 (
            .O(N__25941),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__3859 (
            .O(N__25936),
            .I(N__25933));
    InMux I__3858 (
            .O(N__25933),
            .I(N__25926));
    InMux I__3857 (
            .O(N__25932),
            .I(N__25926));
    InMux I__3856 (
            .O(N__25931),
            .I(N__25923));
    LocalMux I__3855 (
            .O(N__25926),
            .I(N__25920));
    LocalMux I__3854 (
            .O(N__25923),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__3853 (
            .O(N__25920),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__3852 (
            .O(N__25915),
            .I(N__25912));
    LocalMux I__3851 (
            .O(N__25912),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    CascadeMux I__3850 (
            .O(N__25909),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_));
    CascadeMux I__3849 (
            .O(N__25906),
            .I(N__25903));
    InMux I__3848 (
            .O(N__25903),
            .I(N__25897));
    InMux I__3847 (
            .O(N__25902),
            .I(N__25897));
    LocalMux I__3846 (
            .O(N__25897),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    CascadeMux I__3845 (
            .O(N__25894),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__3844 (
            .O(N__25891),
            .I(N__25885));
    InMux I__3843 (
            .O(N__25890),
            .I(N__25885));
    LocalMux I__3842 (
            .O(N__25885),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    CascadeMux I__3841 (
            .O(N__25882),
            .I(N__25879));
    InMux I__3840 (
            .O(N__25879),
            .I(N__25876));
    LocalMux I__3839 (
            .O(N__25876),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__3838 (
            .O(N__25873),
            .I(N__25869));
    InMux I__3837 (
            .O(N__25872),
            .I(N__25866));
    LocalMux I__3836 (
            .O(N__25869),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__3835 (
            .O(N__25866),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__3834 (
            .O(N__25861),
            .I(N__25857));
    InMux I__3833 (
            .O(N__25860),
            .I(N__25854));
    LocalMux I__3832 (
            .O(N__25857),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__3831 (
            .O(N__25854),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__3830 (
            .O(N__25849),
            .I(N__25845));
    CascadeMux I__3829 (
            .O(N__25848),
            .I(N__25842));
    InMux I__3828 (
            .O(N__25845),
            .I(N__25839));
    InMux I__3827 (
            .O(N__25842),
            .I(N__25835));
    LocalMux I__3826 (
            .O(N__25839),
            .I(N__25832));
    InMux I__3825 (
            .O(N__25838),
            .I(N__25829));
    LocalMux I__3824 (
            .O(N__25835),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3823 (
            .O(N__25832),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3822 (
            .O(N__25829),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__3821 (
            .O(N__25822),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    InMux I__3820 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__3819 (
            .O(N__25816),
            .I(N__25813));
    Span12Mux_s11_h I__3818 (
            .O(N__25813),
            .I(N__25810));
    Odrv12 I__3817 (
            .O(N__25810),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    InMux I__3816 (
            .O(N__25807),
            .I(N__25804));
    LocalMux I__3815 (
            .O(N__25804),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    CascadeMux I__3814 (
            .O(N__25801),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    CascadeMux I__3813 (
            .O(N__25798),
            .I(N__25795));
    InMux I__3812 (
            .O(N__25795),
            .I(N__25792));
    LocalMux I__3811 (
            .O(N__25792),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__3810 (
            .O(N__25789),
            .I(N__25786));
    LocalMux I__3809 (
            .O(N__25786),
            .I(N__25783));
    Span4Mux_v I__3808 (
            .O(N__25783),
            .I(N__25780));
    Odrv4 I__3807 (
            .O(N__25780),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__3806 (
            .O(N__25777),
            .I(N__25774));
    LocalMux I__3805 (
            .O(N__25774),
            .I(N__25771));
    Odrv12 I__3804 (
            .O(N__25771),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__3803 (
            .O(N__25768),
            .I(N__25765));
    LocalMux I__3802 (
            .O(N__25765),
            .I(N__25762));
    Odrv12 I__3801 (
            .O(N__25762),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__3800 (
            .O(N__25759),
            .I(N__25755));
    InMux I__3799 (
            .O(N__25758),
            .I(N__25752));
    LocalMux I__3798 (
            .O(N__25755),
            .I(N__25749));
    LocalMux I__3797 (
            .O(N__25752),
            .I(N__25746));
    Span4Mux_h I__3796 (
            .O(N__25749),
            .I(N__25739));
    Span4Mux_v I__3795 (
            .O(N__25746),
            .I(N__25739));
    InMux I__3794 (
            .O(N__25745),
            .I(N__25734));
    InMux I__3793 (
            .O(N__25744),
            .I(N__25734));
    Odrv4 I__3792 (
            .O(N__25739),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__3791 (
            .O(N__25734),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    CascadeMux I__3790 (
            .O(N__25729),
            .I(N__25726));
    InMux I__3789 (
            .O(N__25726),
            .I(N__25723));
    LocalMux I__3788 (
            .O(N__25723),
            .I(N__25720));
    Span12Mux_h I__3787 (
            .O(N__25720),
            .I(N__25717));
    Odrv12 I__3786 (
            .O(N__25717),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__3785 (
            .O(N__25714),
            .I(N__25711));
    InMux I__3784 (
            .O(N__25711),
            .I(N__25708));
    LocalMux I__3783 (
            .O(N__25708),
            .I(N__25705));
    Span4Mux_v I__3782 (
            .O(N__25705),
            .I(N__25702));
    Span4Mux_v I__3781 (
            .O(N__25702),
            .I(N__25699));
    Odrv4 I__3780 (
            .O(N__25699),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__3779 (
            .O(N__25696),
            .I(N__25693));
    InMux I__3778 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__3777 (
            .O(N__25690),
            .I(N__25687));
    Sp12to4 I__3776 (
            .O(N__25687),
            .I(N__25684));
    Odrv12 I__3775 (
            .O(N__25684),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    CascadeMux I__3774 (
            .O(N__25681),
            .I(N__25678));
    InMux I__3773 (
            .O(N__25678),
            .I(N__25675));
    LocalMux I__3772 (
            .O(N__25675),
            .I(N__25672));
    Span4Mux_v I__3771 (
            .O(N__25672),
            .I(N__25669));
    Span4Mux_h I__3770 (
            .O(N__25669),
            .I(N__25666));
    Odrv4 I__3769 (
            .O(N__25666),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    CascadeMux I__3768 (
            .O(N__25663),
            .I(N__25660));
    InMux I__3767 (
            .O(N__25660),
            .I(N__25657));
    LocalMux I__3766 (
            .O(N__25657),
            .I(N__25654));
    Span4Mux_v I__3765 (
            .O(N__25654),
            .I(N__25651));
    Span4Mux_v I__3764 (
            .O(N__25651),
            .I(N__25648));
    Odrv4 I__3763 (
            .O(N__25648),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__3762 (
            .O(N__25645),
            .I(N__25642));
    InMux I__3761 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__3760 (
            .O(N__25639),
            .I(N__25636));
    Span4Mux_v I__3759 (
            .O(N__25636),
            .I(N__25633));
    Odrv4 I__3758 (
            .O(N__25633),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__3757 (
            .O(N__25630),
            .I(N__25624));
    InMux I__3756 (
            .O(N__25629),
            .I(N__25624));
    LocalMux I__3755 (
            .O(N__25624),
            .I(N__25619));
    InMux I__3754 (
            .O(N__25623),
            .I(N__25614));
    InMux I__3753 (
            .O(N__25622),
            .I(N__25614));
    Odrv4 I__3752 (
            .O(N__25619),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__3751 (
            .O(N__25614),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__3750 (
            .O(N__25609),
            .I(N__25606));
    LocalMux I__3749 (
            .O(N__25606),
            .I(N__25603));
    Odrv12 I__3748 (
            .O(N__25603),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__3747 (
            .O(N__25600),
            .I(N__25597));
    LocalMux I__3746 (
            .O(N__25597),
            .I(N__25594));
    Span4Mux_v I__3745 (
            .O(N__25594),
            .I(N__25591));
    Odrv4 I__3744 (
            .O(N__25591),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__3743 (
            .O(N__25588),
            .I(N__25585));
    LocalMux I__3742 (
            .O(N__25585),
            .I(N__25582));
    Span4Mux_v I__3741 (
            .O(N__25582),
            .I(N__25579));
    Odrv4 I__3740 (
            .O(N__25579),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__3739 (
            .O(N__25576),
            .I(N__25573));
    InMux I__3738 (
            .O(N__25573),
            .I(N__25570));
    LocalMux I__3737 (
            .O(N__25570),
            .I(N__25567));
    Span4Mux_v I__3736 (
            .O(N__25567),
            .I(N__25564));
    Odrv4 I__3735 (
            .O(N__25564),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__3734 (
            .O(N__25561),
            .I(N__25558));
    LocalMux I__3733 (
            .O(N__25558),
            .I(N__25555));
    Span4Mux_v I__3732 (
            .O(N__25555),
            .I(N__25552));
    Odrv4 I__3731 (
            .O(N__25552),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__3730 (
            .O(N__25549),
            .I(N__25546));
    LocalMux I__3729 (
            .O(N__25546),
            .I(N__25543));
    Span4Mux_v I__3728 (
            .O(N__25543),
            .I(N__25540));
    Odrv4 I__3727 (
            .O(N__25540),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__3726 (
            .O(N__25537),
            .I(N__25534));
    LocalMux I__3725 (
            .O(N__25534),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__3724 (
            .O(N__25531),
            .I(N__25528));
    InMux I__3723 (
            .O(N__25528),
            .I(N__25525));
    LocalMux I__3722 (
            .O(N__25525),
            .I(N__25522));
    Span4Mux_v I__3721 (
            .O(N__25522),
            .I(N__25519));
    Odrv4 I__3720 (
            .O(N__25519),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    InMux I__3719 (
            .O(N__25516),
            .I(N__25513));
    LocalMux I__3718 (
            .O(N__25513),
            .I(N__25510));
    Odrv4 I__3717 (
            .O(N__25510),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__3716 (
            .O(N__25507),
            .I(N__25504));
    LocalMux I__3715 (
            .O(N__25504),
            .I(N__25501));
    Odrv4 I__3714 (
            .O(N__25501),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__3713 (
            .O(N__25498),
            .I(N__25495));
    LocalMux I__3712 (
            .O(N__25495),
            .I(N__25492));
    Span4Mux_v I__3711 (
            .O(N__25492),
            .I(N__25489));
    Odrv4 I__3710 (
            .O(N__25489),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__3709 (
            .O(N__25486),
            .I(N__25483));
    InMux I__3708 (
            .O(N__25483),
            .I(N__25480));
    LocalMux I__3707 (
            .O(N__25480),
            .I(N__25477));
    Span4Mux_v I__3706 (
            .O(N__25477),
            .I(N__25474));
    Odrv4 I__3705 (
            .O(N__25474),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    CascadeMux I__3704 (
            .O(N__25471),
            .I(N__25468));
    InMux I__3703 (
            .O(N__25468),
            .I(N__25465));
    LocalMux I__3702 (
            .O(N__25465),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__3701 (
            .O(N__25462),
            .I(N__25459));
    InMux I__3700 (
            .O(N__25459),
            .I(N__25456));
    LocalMux I__3699 (
            .O(N__25456),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__3698 (
            .O(N__25453),
            .I(N__25450));
    InMux I__3697 (
            .O(N__25450),
            .I(N__25447));
    LocalMux I__3696 (
            .O(N__25447),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    CascadeMux I__3695 (
            .O(N__25444),
            .I(N__25441));
    InMux I__3694 (
            .O(N__25441),
            .I(N__25438));
    LocalMux I__3693 (
            .O(N__25438),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__3692 (
            .O(N__25435),
            .I(N__25432));
    LocalMux I__3691 (
            .O(N__25432),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__3690 (
            .O(N__25429),
            .I(N__25426));
    InMux I__3689 (
            .O(N__25426),
            .I(N__25423));
    LocalMux I__3688 (
            .O(N__25423),
            .I(N__25420));
    Span4Mux_v I__3687 (
            .O(N__25420),
            .I(N__25417));
    Odrv4 I__3686 (
            .O(N__25417),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__3685 (
            .O(N__25414),
            .I(N__25411));
    LocalMux I__3684 (
            .O(N__25411),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__3683 (
            .O(N__25408),
            .I(N__25405));
    InMux I__3682 (
            .O(N__25405),
            .I(N__25402));
    LocalMux I__3681 (
            .O(N__25402),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__3680 (
            .O(N__25399),
            .I(N__25396));
    LocalMux I__3679 (
            .O(N__25396),
            .I(N__25393));
    Odrv12 I__3678 (
            .O(N__25393),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__3677 (
            .O(N__25390),
            .I(N__25387));
    LocalMux I__3676 (
            .O(N__25387),
            .I(N__25384));
    Odrv12 I__3675 (
            .O(N__25384),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__3674 (
            .O(N__25381),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    CascadeMux I__3673 (
            .O(N__25378),
            .I(N__25353));
    InMux I__3672 (
            .O(N__25377),
            .I(N__25342));
    InMux I__3671 (
            .O(N__25376),
            .I(N__25342));
    InMux I__3670 (
            .O(N__25375),
            .I(N__25327));
    InMux I__3669 (
            .O(N__25374),
            .I(N__25327));
    InMux I__3668 (
            .O(N__25373),
            .I(N__25327));
    InMux I__3667 (
            .O(N__25372),
            .I(N__25327));
    InMux I__3666 (
            .O(N__25371),
            .I(N__25327));
    InMux I__3665 (
            .O(N__25370),
            .I(N__25327));
    InMux I__3664 (
            .O(N__25369),
            .I(N__25327));
    InMux I__3663 (
            .O(N__25368),
            .I(N__25310));
    InMux I__3662 (
            .O(N__25367),
            .I(N__25310));
    InMux I__3661 (
            .O(N__25366),
            .I(N__25310));
    InMux I__3660 (
            .O(N__25365),
            .I(N__25310));
    InMux I__3659 (
            .O(N__25364),
            .I(N__25310));
    InMux I__3658 (
            .O(N__25363),
            .I(N__25310));
    InMux I__3657 (
            .O(N__25362),
            .I(N__25310));
    InMux I__3656 (
            .O(N__25361),
            .I(N__25310));
    InMux I__3655 (
            .O(N__25360),
            .I(N__25299));
    InMux I__3654 (
            .O(N__25359),
            .I(N__25299));
    InMux I__3653 (
            .O(N__25358),
            .I(N__25299));
    InMux I__3652 (
            .O(N__25357),
            .I(N__25299));
    InMux I__3651 (
            .O(N__25356),
            .I(N__25299));
    InMux I__3650 (
            .O(N__25353),
            .I(N__25296));
    InMux I__3649 (
            .O(N__25352),
            .I(N__25280));
    InMux I__3648 (
            .O(N__25351),
            .I(N__25280));
    InMux I__3647 (
            .O(N__25350),
            .I(N__25280));
    InMux I__3646 (
            .O(N__25349),
            .I(N__25280));
    InMux I__3645 (
            .O(N__25348),
            .I(N__25280));
    InMux I__3644 (
            .O(N__25347),
            .I(N__25280));
    LocalMux I__3643 (
            .O(N__25342),
            .I(N__25271));
    LocalMux I__3642 (
            .O(N__25327),
            .I(N__25271));
    LocalMux I__3641 (
            .O(N__25310),
            .I(N__25271));
    LocalMux I__3640 (
            .O(N__25299),
            .I(N__25271));
    LocalMux I__3639 (
            .O(N__25296),
            .I(N__25268));
    InMux I__3638 (
            .O(N__25295),
            .I(N__25263));
    InMux I__3637 (
            .O(N__25294),
            .I(N__25263));
    InMux I__3636 (
            .O(N__25293),
            .I(N__25260));
    LocalMux I__3635 (
            .O(N__25280),
            .I(N__25255));
    Span4Mux_v I__3634 (
            .O(N__25271),
            .I(N__25255));
    Odrv4 I__3633 (
            .O(N__25268),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__3632 (
            .O(N__25263),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__3631 (
            .O(N__25260),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__3630 (
            .O(N__25255),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__3629 (
            .O(N__25246),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__3628 (
            .O(N__25243),
            .I(N__25240));
    LocalMux I__3627 (
            .O(N__25240),
            .I(N__25237));
    Span4Mux_h I__3626 (
            .O(N__25237),
            .I(N__25234));
    Odrv4 I__3625 (
            .O(N__25234),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__3624 (
            .O(N__25231),
            .I(N__25228));
    LocalMux I__3623 (
            .O(N__25228),
            .I(N__25225));
    Odrv4 I__3622 (
            .O(N__25225),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__3621 (
            .O(N__25222),
            .I(N__25219));
    LocalMux I__3620 (
            .O(N__25219),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__3619 (
            .O(N__25216),
            .I(N__25213));
    InMux I__3618 (
            .O(N__25213),
            .I(N__25210));
    LocalMux I__3617 (
            .O(N__25210),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    CascadeMux I__3616 (
            .O(N__25207),
            .I(N__25204));
    InMux I__3615 (
            .O(N__25204),
            .I(N__25201));
    LocalMux I__3614 (
            .O(N__25201),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    CascadeMux I__3613 (
            .O(N__25198),
            .I(N__25195));
    InMux I__3612 (
            .O(N__25195),
            .I(N__25192));
    LocalMux I__3611 (
            .O(N__25192),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__3610 (
            .O(N__25189),
            .I(N__25186));
    LocalMux I__3609 (
            .O(N__25186),
            .I(N__25183));
    Odrv4 I__3608 (
            .O(N__25183),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__3607 (
            .O(N__25180),
            .I(N__25177));
    LocalMux I__3606 (
            .O(N__25177),
            .I(N__25174));
    Span4Mux_h I__3605 (
            .O(N__25174),
            .I(N__25171));
    Odrv4 I__3604 (
            .O(N__25171),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__3603 (
            .O(N__25168),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__3602 (
            .O(N__25165),
            .I(N__25162));
    LocalMux I__3601 (
            .O(N__25162),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__3600 (
            .O(N__25159),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__3599 (
            .O(N__25156),
            .I(N__25153));
    LocalMux I__3598 (
            .O(N__25153),
            .I(N__25150));
    Odrv4 I__3597 (
            .O(N__25150),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__3596 (
            .O(N__25147),
            .I(bfn_10_17_0_));
    InMux I__3595 (
            .O(N__25144),
            .I(N__25141));
    LocalMux I__3594 (
            .O(N__25141),
            .I(N__25138));
    Odrv12 I__3593 (
            .O(N__25138),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__3592 (
            .O(N__25135),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__3591 (
            .O(N__25132),
            .I(N__25129));
    LocalMux I__3590 (
            .O(N__25129),
            .I(N__25126));
    Odrv4 I__3589 (
            .O(N__25126),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__3588 (
            .O(N__25123),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__3587 (
            .O(N__25120),
            .I(N__25117));
    LocalMux I__3586 (
            .O(N__25117),
            .I(N__25114));
    Odrv12 I__3585 (
            .O(N__25114),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__3584 (
            .O(N__25111),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__3583 (
            .O(N__25108),
            .I(N__25105));
    LocalMux I__3582 (
            .O(N__25105),
            .I(N__25102));
    Span4Mux_h I__3581 (
            .O(N__25102),
            .I(N__25099));
    Odrv4 I__3580 (
            .O(N__25099),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__3579 (
            .O(N__25096),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__3578 (
            .O(N__25093),
            .I(N__25090));
    LocalMux I__3577 (
            .O(N__25090),
            .I(N__25087));
    Odrv4 I__3576 (
            .O(N__25087),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__3575 (
            .O(N__25084),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__3574 (
            .O(N__25081),
            .I(N__25078));
    LocalMux I__3573 (
            .O(N__25078),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__3572 (
            .O(N__25075),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__3571 (
            .O(N__25072),
            .I(N__25069));
    LocalMux I__3570 (
            .O(N__25069),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__3569 (
            .O(N__25066),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__3568 (
            .O(N__25063),
            .I(N__25060));
    LocalMux I__3567 (
            .O(N__25060),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__3566 (
            .O(N__25057),
            .I(bfn_10_16_0_));
    InMux I__3565 (
            .O(N__25054),
            .I(N__25051));
    LocalMux I__3564 (
            .O(N__25051),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__3563 (
            .O(N__25048),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__3562 (
            .O(N__25045),
            .I(N__25042));
    LocalMux I__3561 (
            .O(N__25042),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__3560 (
            .O(N__25039),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__3559 (
            .O(N__25036),
            .I(N__25033));
    LocalMux I__3558 (
            .O(N__25033),
            .I(N__25030));
    Odrv4 I__3557 (
            .O(N__25030),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__3556 (
            .O(N__25027),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__3555 (
            .O(N__25024),
            .I(N__25021));
    LocalMux I__3554 (
            .O(N__25021),
            .I(N__25018));
    Span4Mux_h I__3553 (
            .O(N__25018),
            .I(N__25015));
    Odrv4 I__3552 (
            .O(N__25015),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__3551 (
            .O(N__25012),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__3550 (
            .O(N__25009),
            .I(N__25006));
    LocalMux I__3549 (
            .O(N__25006),
            .I(N__25003));
    Odrv4 I__3548 (
            .O(N__25003),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__3547 (
            .O(N__25000),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__3546 (
            .O(N__24997),
            .I(N__24994));
    LocalMux I__3545 (
            .O(N__24994),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__3544 (
            .O(N__24991),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__3543 (
            .O(N__24988),
            .I(N__24985));
    LocalMux I__3542 (
            .O(N__24985),
            .I(N__24982));
    Odrv4 I__3541 (
            .O(N__24982),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__3540 (
            .O(N__24979),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__3539 (
            .O(N__24976),
            .I(N__24973));
    LocalMux I__3538 (
            .O(N__24973),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__3537 (
            .O(N__24970),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__3536 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__3535 (
            .O(N__24964),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__3534 (
            .O(N__24961),
            .I(bfn_10_15_0_));
    InMux I__3533 (
            .O(N__24958),
            .I(N__24955));
    LocalMux I__3532 (
            .O(N__24955),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__3531 (
            .O(N__24952),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__3530 (
            .O(N__24949),
            .I(N__24946));
    LocalMux I__3529 (
            .O(N__24946),
            .I(N__24943));
    Span4Mux_v I__3528 (
            .O(N__24943),
            .I(N__24940));
    Odrv4 I__3527 (
            .O(N__24940),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__3526 (
            .O(N__24937),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__3525 (
            .O(N__24934),
            .I(N__24931));
    LocalMux I__3524 (
            .O(N__24931),
            .I(N__24928));
    Odrv4 I__3523 (
            .O(N__24928),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__3522 (
            .O(N__24925),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__3521 (
            .O(N__24922),
            .I(N__24919));
    LocalMux I__3520 (
            .O(N__24919),
            .I(N__24916));
    Odrv4 I__3519 (
            .O(N__24916),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__3518 (
            .O(N__24913),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__3517 (
            .O(N__24910),
            .I(N__24907));
    LocalMux I__3516 (
            .O(N__24907),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__3515 (
            .O(N__24904),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__3514 (
            .O(N__24901),
            .I(N__24896));
    InMux I__3513 (
            .O(N__24900),
            .I(N__24893));
    InMux I__3512 (
            .O(N__24899),
            .I(N__24890));
    LocalMux I__3511 (
            .O(N__24896),
            .I(N__24887));
    LocalMux I__3510 (
            .O(N__24893),
            .I(N__24884));
    LocalMux I__3509 (
            .O(N__24890),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv12 I__3508 (
            .O(N__24887),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__3507 (
            .O(N__24884),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__3506 (
            .O(N__24877),
            .I(N__24872));
    InMux I__3505 (
            .O(N__24876),
            .I(N__24869));
    InMux I__3504 (
            .O(N__24875),
            .I(N__24866));
    LocalMux I__3503 (
            .O(N__24872),
            .I(N__24863));
    LocalMux I__3502 (
            .O(N__24869),
            .I(N__24860));
    LocalMux I__3501 (
            .O(N__24866),
            .I(N__24857));
    Span4Mux_v I__3500 (
            .O(N__24863),
            .I(N__24853));
    Span4Mux_v I__3499 (
            .O(N__24860),
            .I(N__24848));
    Span4Mux_v I__3498 (
            .O(N__24857),
            .I(N__24848));
    InMux I__3497 (
            .O(N__24856),
            .I(N__24845));
    Odrv4 I__3496 (
            .O(N__24853),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__3495 (
            .O(N__24848),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__3494 (
            .O(N__24845),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__3493 (
            .O(N__24838),
            .I(N__24833));
    InMux I__3492 (
            .O(N__24837),
            .I(N__24828));
    InMux I__3491 (
            .O(N__24836),
            .I(N__24828));
    LocalMux I__3490 (
            .O(N__24833),
            .I(N__24824));
    LocalMux I__3489 (
            .O(N__24828),
            .I(N__24821));
    InMux I__3488 (
            .O(N__24827),
            .I(N__24818));
    Span4Mux_v I__3487 (
            .O(N__24824),
            .I(N__24813));
    Span4Mux_v I__3486 (
            .O(N__24821),
            .I(N__24813));
    LocalMux I__3485 (
            .O(N__24818),
            .I(N__24810));
    Odrv4 I__3484 (
            .O(N__24813),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__3483 (
            .O(N__24810),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__3482 (
            .O(N__24805),
            .I(N__24802));
    LocalMux I__3481 (
            .O(N__24802),
            .I(N__24798));
    InMux I__3480 (
            .O(N__24801),
            .I(N__24795));
    Odrv4 I__3479 (
            .O(N__24798),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    LocalMux I__3478 (
            .O(N__24795),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__3477 (
            .O(N__24790),
            .I(N__24787));
    LocalMux I__3476 (
            .O(N__24787),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__3475 (
            .O(N__24784),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__3474 (
            .O(N__24781),
            .I(N__24778));
    LocalMux I__3473 (
            .O(N__24778),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__3472 (
            .O(N__24775),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    CascadeMux I__3471 (
            .O(N__24772),
            .I(elapsed_time_ns_1_RNI58DN9_0_27_cascade_));
    CascadeMux I__3470 (
            .O(N__24769),
            .I(N__24765));
    InMux I__3469 (
            .O(N__24768),
            .I(N__24760));
    InMux I__3468 (
            .O(N__24765),
            .I(N__24760));
    LocalMux I__3467 (
            .O(N__24760),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    CascadeMux I__3466 (
            .O(N__24757),
            .I(elapsed_time_ns_1_RNI47DN9_0_26_cascade_));
    InMux I__3465 (
            .O(N__24754),
            .I(N__24748));
    InMux I__3464 (
            .O(N__24753),
            .I(N__24748));
    LocalMux I__3463 (
            .O(N__24748),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    CascadeMux I__3462 (
            .O(N__24745),
            .I(N__24742));
    InMux I__3461 (
            .O(N__24742),
            .I(N__24739));
    LocalMux I__3460 (
            .O(N__24739),
            .I(N__24736));
    Span4Mux_h I__3459 (
            .O(N__24736),
            .I(N__24733));
    Odrv4 I__3458 (
            .O(N__24733),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    CascadeMux I__3457 (
            .O(N__24730),
            .I(N__24726));
    InMux I__3456 (
            .O(N__24729),
            .I(N__24721));
    InMux I__3455 (
            .O(N__24726),
            .I(N__24721));
    LocalMux I__3454 (
            .O(N__24721),
            .I(N__24718));
    Odrv12 I__3453 (
            .O(N__24718),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__3452 (
            .O(N__24715),
            .I(N__24711));
    InMux I__3451 (
            .O(N__24714),
            .I(N__24705));
    InMux I__3450 (
            .O(N__24711),
            .I(N__24705));
    InMux I__3449 (
            .O(N__24710),
            .I(N__24702));
    LocalMux I__3448 (
            .O(N__24705),
            .I(N__24699));
    LocalMux I__3447 (
            .O(N__24702),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__3446 (
            .O(N__24699),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__3445 (
            .O(N__24694),
            .I(N__24687));
    InMux I__3444 (
            .O(N__24693),
            .I(N__24687));
    InMux I__3443 (
            .O(N__24692),
            .I(N__24684));
    LocalMux I__3442 (
            .O(N__24687),
            .I(N__24681));
    LocalMux I__3441 (
            .O(N__24684),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__3440 (
            .O(N__24681),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__3439 (
            .O(N__24676),
            .I(N__24673));
    LocalMux I__3438 (
            .O(N__24673),
            .I(N__24670));
    Odrv4 I__3437 (
            .O(N__24670),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    CascadeMux I__3436 (
            .O(N__24667),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__3435 (
            .O(N__24664),
            .I(N__24658));
    InMux I__3434 (
            .O(N__24663),
            .I(N__24658));
    LocalMux I__3433 (
            .O(N__24658),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    CascadeMux I__3432 (
            .O(N__24655),
            .I(N__24652));
    InMux I__3431 (
            .O(N__24652),
            .I(N__24649));
    LocalMux I__3430 (
            .O(N__24649),
            .I(N__24646));
    Odrv12 I__3429 (
            .O(N__24646),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__3428 (
            .O(N__24643),
            .I(N__24640));
    LocalMux I__3427 (
            .O(N__24640),
            .I(N__24637));
    Span4Mux_h I__3426 (
            .O(N__24637),
            .I(N__24634));
    Odrv4 I__3425 (
            .O(N__24634),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__3424 (
            .O(N__24631),
            .I(N__24628));
    InMux I__3423 (
            .O(N__24628),
            .I(N__24625));
    LocalMux I__3422 (
            .O(N__24625),
            .I(N__24622));
    Odrv12 I__3421 (
            .O(N__24622),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__3420 (
            .O(N__24619),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__3419 (
            .O(N__24616),
            .I(N__24613));
    InMux I__3418 (
            .O(N__24613),
            .I(N__24610));
    LocalMux I__3417 (
            .O(N__24610),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    CascadeMux I__3416 (
            .O(N__24607),
            .I(elapsed_time_ns_1_RNII43T9_0_6_cascade_));
    CascadeMux I__3415 (
            .O(N__24604),
            .I(N__24601));
    InMux I__3414 (
            .O(N__24601),
            .I(N__24598));
    LocalMux I__3413 (
            .O(N__24598),
            .I(N__24595));
    Odrv4 I__3412 (
            .O(N__24595),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__3411 (
            .O(N__24592),
            .I(N__24587));
    InMux I__3410 (
            .O(N__24591),
            .I(N__24584));
    InMux I__3409 (
            .O(N__24590),
            .I(N__24579));
    InMux I__3408 (
            .O(N__24587),
            .I(N__24579));
    LocalMux I__3407 (
            .O(N__24584),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__3406 (
            .O(N__24579),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__3405 (
            .O(N__24574),
            .I(N__24569));
    InMux I__3404 (
            .O(N__24573),
            .I(N__24564));
    InMux I__3403 (
            .O(N__24572),
            .I(N__24564));
    LocalMux I__3402 (
            .O(N__24569),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__3401 (
            .O(N__24564),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__3400 (
            .O(N__24559),
            .I(N__24556));
    LocalMux I__3399 (
            .O(N__24556),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__3398 (
            .O(N__24553),
            .I(N__24550));
    LocalMux I__3397 (
            .O(N__24550),
            .I(N__24547));
    Span4Mux_h I__3396 (
            .O(N__24547),
            .I(N__24544));
    Span4Mux_h I__3395 (
            .O(N__24544),
            .I(N__24541));
    Odrv4 I__3394 (
            .O(N__24541),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__3393 (
            .O(N__24538),
            .I(N__24534));
    InMux I__3392 (
            .O(N__24537),
            .I(N__24531));
    LocalMux I__3391 (
            .O(N__24534),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3390 (
            .O(N__24531),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__3389 (
            .O(N__24526),
            .I(N__24523));
    InMux I__3388 (
            .O(N__24523),
            .I(N__24520));
    LocalMux I__3387 (
            .O(N__24520),
            .I(N__24517));
    Odrv4 I__3386 (
            .O(N__24517),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__3385 (
            .O(N__24514),
            .I(N__24511));
    LocalMux I__3384 (
            .O(N__24511),
            .I(N__24508));
    Span4Mux_h I__3383 (
            .O(N__24508),
            .I(N__24505));
    Odrv4 I__3382 (
            .O(N__24505),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__3381 (
            .O(N__24502),
            .I(N__24498));
    InMux I__3380 (
            .O(N__24501),
            .I(N__24495));
    LocalMux I__3379 (
            .O(N__24498),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3378 (
            .O(N__24495),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__3377 (
            .O(N__24490),
            .I(N__24487));
    InMux I__3376 (
            .O(N__24487),
            .I(N__24484));
    LocalMux I__3375 (
            .O(N__24484),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__3374 (
            .O(N__24481),
            .I(N__24478));
    LocalMux I__3373 (
            .O(N__24478),
            .I(N__24475));
    Odrv4 I__3372 (
            .O(N__24475),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__3371 (
            .O(N__24472),
            .I(N__24468));
    InMux I__3370 (
            .O(N__24471),
            .I(N__24465));
    LocalMux I__3369 (
            .O(N__24468),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3368 (
            .O(N__24465),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__3367 (
            .O(N__24460),
            .I(N__24457));
    InMux I__3366 (
            .O(N__24457),
            .I(N__24454));
    LocalMux I__3365 (
            .O(N__24454),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3364 (
            .O(N__24451),
            .I(N__24448));
    LocalMux I__3363 (
            .O(N__24448),
            .I(N__24445));
    Span4Mux_h I__3362 (
            .O(N__24445),
            .I(N__24442));
    Odrv4 I__3361 (
            .O(N__24442),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    CascadeMux I__3360 (
            .O(N__24439),
            .I(N__24436));
    InMux I__3359 (
            .O(N__24436),
            .I(N__24433));
    LocalMux I__3358 (
            .O(N__24433),
            .I(N__24430));
    Span4Mux_h I__3357 (
            .O(N__24430),
            .I(N__24427));
    Odrv4 I__3356 (
            .O(N__24427),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__3355 (
            .O(N__24424),
            .I(N__24421));
    LocalMux I__3354 (
            .O(N__24421),
            .I(N__24418));
    Span4Mux_h I__3353 (
            .O(N__24418),
            .I(N__24415));
    Odrv4 I__3352 (
            .O(N__24415),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__3351 (
            .O(N__24412),
            .I(N__24409));
    InMux I__3350 (
            .O(N__24409),
            .I(N__24406));
    LocalMux I__3349 (
            .O(N__24406),
            .I(N__24403));
    Span4Mux_h I__3348 (
            .O(N__24403),
            .I(N__24400));
    Odrv4 I__3347 (
            .O(N__24400),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__3346 (
            .O(N__24397),
            .I(N__24394));
    LocalMux I__3345 (
            .O(N__24394),
            .I(N__24391));
    Odrv4 I__3344 (
            .O(N__24391),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    CascadeMux I__3343 (
            .O(N__24388),
            .I(N__24385));
    InMux I__3342 (
            .O(N__24385),
            .I(N__24382));
    LocalMux I__3341 (
            .O(N__24382),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__3340 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__3339 (
            .O(N__24376),
            .I(N__24373));
    Odrv4 I__3338 (
            .O(N__24373),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__3337 (
            .O(N__24370),
            .I(N__24366));
    InMux I__3336 (
            .O(N__24369),
            .I(N__24363));
    LocalMux I__3335 (
            .O(N__24366),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3334 (
            .O(N__24363),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__3333 (
            .O(N__24358),
            .I(N__24355));
    InMux I__3332 (
            .O(N__24355),
            .I(N__24352));
    LocalMux I__3331 (
            .O(N__24352),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3330 (
            .O(N__24349),
            .I(N__24345));
    InMux I__3329 (
            .O(N__24348),
            .I(N__24342));
    LocalMux I__3328 (
            .O(N__24345),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3327 (
            .O(N__24342),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3326 (
            .O(N__24337),
            .I(N__24334));
    LocalMux I__3325 (
            .O(N__24334),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3324 (
            .O(N__24331),
            .I(N__24327));
    InMux I__3323 (
            .O(N__24330),
            .I(N__24324));
    LocalMux I__3322 (
            .O(N__24327),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3321 (
            .O(N__24324),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__3320 (
            .O(N__24319),
            .I(N__24316));
    InMux I__3319 (
            .O(N__24316),
            .I(N__24313));
    LocalMux I__3318 (
            .O(N__24313),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__3317 (
            .O(N__24310),
            .I(N__24306));
    InMux I__3316 (
            .O(N__24309),
            .I(N__24303));
    LocalMux I__3315 (
            .O(N__24306),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__3314 (
            .O(N__24303),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3313 (
            .O(N__24298),
            .I(N__24295));
    LocalMux I__3312 (
            .O(N__24295),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3311 (
            .O(N__24292),
            .I(N__24288));
    InMux I__3310 (
            .O(N__24291),
            .I(N__24285));
    LocalMux I__3309 (
            .O(N__24288),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3308 (
            .O(N__24285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3307 (
            .O(N__24280),
            .I(N__24277));
    LocalMux I__3306 (
            .O(N__24277),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__3305 (
            .O(N__24274),
            .I(N__24270));
    InMux I__3304 (
            .O(N__24273),
            .I(N__24267));
    LocalMux I__3303 (
            .O(N__24270),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3302 (
            .O(N__24267),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3301 (
            .O(N__24262),
            .I(N__24259));
    LocalMux I__3300 (
            .O(N__24259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__3299 (
            .O(N__24256),
            .I(N__24252));
    InMux I__3298 (
            .O(N__24255),
            .I(N__24249));
    LocalMux I__3297 (
            .O(N__24252),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3296 (
            .O(N__24249),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__3295 (
            .O(N__24244),
            .I(N__24241));
    InMux I__3294 (
            .O(N__24241),
            .I(N__24238));
    LocalMux I__3293 (
            .O(N__24238),
            .I(N__24235));
    Odrv4 I__3292 (
            .O(N__24235),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__3291 (
            .O(N__24232),
            .I(N__24228));
    InMux I__3290 (
            .O(N__24231),
            .I(N__24225));
    LocalMux I__3289 (
            .O(N__24228),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3288 (
            .O(N__24225),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__3287 (
            .O(N__24220),
            .I(N__24217));
    InMux I__3286 (
            .O(N__24217),
            .I(N__24214));
    LocalMux I__3285 (
            .O(N__24214),
            .I(N__24211));
    Odrv4 I__3284 (
            .O(N__24211),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__3283 (
            .O(N__24208),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    CascadeMux I__3282 (
            .O(N__24205),
            .I(N__24202));
    InMux I__3281 (
            .O(N__24202),
            .I(N__24199));
    LocalMux I__3280 (
            .O(N__24199),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ));
    CascadeMux I__3279 (
            .O(N__24196),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__3278 (
            .O(N__24193),
            .I(N__24190));
    LocalMux I__3277 (
            .O(N__24190),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__3276 (
            .O(N__24187),
            .I(N__24184));
    LocalMux I__3275 (
            .O(N__24184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__3274 (
            .O(N__24181),
            .I(N__24178));
    LocalMux I__3273 (
            .O(N__24178),
            .I(N__24175));
    Odrv4 I__3272 (
            .O(N__24175),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__3271 (
            .O(N__24172),
            .I(N__24168));
    InMux I__3270 (
            .O(N__24171),
            .I(N__24165));
    LocalMux I__3269 (
            .O(N__24168),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3268 (
            .O(N__24165),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__3267 (
            .O(N__24160),
            .I(N__24157));
    InMux I__3266 (
            .O(N__24157),
            .I(N__24154));
    LocalMux I__3265 (
            .O(N__24154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__3264 (
            .O(N__24151),
            .I(N__24147));
    InMux I__3263 (
            .O(N__24150),
            .I(N__24144));
    LocalMux I__3262 (
            .O(N__24147),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3261 (
            .O(N__24144),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3260 (
            .O(N__24139),
            .I(N__24136));
    LocalMux I__3259 (
            .O(N__24136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__3258 (
            .O(N__24133),
            .I(N__24130));
    LocalMux I__3257 (
            .O(N__24130),
            .I(N__24127));
    Odrv4 I__3256 (
            .O(N__24127),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__3255 (
            .O(N__24124),
            .I(N__24120));
    InMux I__3254 (
            .O(N__24123),
            .I(N__24117));
    LocalMux I__3253 (
            .O(N__24120),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3252 (
            .O(N__24117),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__3251 (
            .O(N__24112),
            .I(N__24109));
    InMux I__3250 (
            .O(N__24109),
            .I(N__24106));
    LocalMux I__3249 (
            .O(N__24106),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__3248 (
            .O(N__24103),
            .I(N__24099));
    InMux I__3247 (
            .O(N__24102),
            .I(N__24096));
    LocalMux I__3246 (
            .O(N__24099),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    LocalMux I__3245 (
            .O(N__24096),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__3244 (
            .O(N__24091),
            .I(N__24087));
    InMux I__3243 (
            .O(N__24090),
            .I(N__24083));
    InMux I__3242 (
            .O(N__24087),
            .I(N__24080));
    InMux I__3241 (
            .O(N__24086),
            .I(N__24077));
    LocalMux I__3240 (
            .O(N__24083),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__3239 (
            .O(N__24080),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__3238 (
            .O(N__24077),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__3237 (
            .O(N__24070),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__3236 (
            .O(N__24067),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    IoInMux I__3235 (
            .O(N__24064),
            .I(N__24061));
    LocalMux I__3234 (
            .O(N__24061),
            .I(N__24058));
    Span4Mux_s1_v I__3233 (
            .O(N__24058),
            .I(N__24055));
    Span4Mux_v I__3232 (
            .O(N__24055),
            .I(N__24051));
    InMux I__3231 (
            .O(N__24054),
            .I(N__24048));
    Sp12to4 I__3230 (
            .O(N__24051),
            .I(N__24044));
    LocalMux I__3229 (
            .O(N__24048),
            .I(N__24041));
    InMux I__3228 (
            .O(N__24047),
            .I(N__24038));
    Odrv12 I__3227 (
            .O(N__24044),
            .I(s1_phy_c));
    Odrv4 I__3226 (
            .O(N__24041),
            .I(s1_phy_c));
    LocalMux I__3225 (
            .O(N__24038),
            .I(s1_phy_c));
    InMux I__3224 (
            .O(N__24031),
            .I(N__24026));
    InMux I__3223 (
            .O(N__24030),
            .I(N__24021));
    InMux I__3222 (
            .O(N__24029),
            .I(N__24021));
    LocalMux I__3221 (
            .O(N__24026),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    LocalMux I__3220 (
            .O(N__24021),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__3219 (
            .O(N__24016),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__3218 (
            .O(N__24013),
            .I(N__24009));
    InMux I__3217 (
            .O(N__24012),
            .I(N__24005));
    InMux I__3216 (
            .O(N__24009),
            .I(N__24002));
    InMux I__3215 (
            .O(N__24008),
            .I(N__23999));
    LocalMux I__3214 (
            .O(N__24005),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__3213 (
            .O(N__24002),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__3212 (
            .O(N__23999),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__3211 (
            .O(N__23992),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__3210 (
            .O(N__23989),
            .I(N__23984));
    CascadeMux I__3209 (
            .O(N__23988),
            .I(N__23981));
    InMux I__3208 (
            .O(N__23987),
            .I(N__23978));
    InMux I__3207 (
            .O(N__23984),
            .I(N__23973));
    InMux I__3206 (
            .O(N__23981),
            .I(N__23973));
    LocalMux I__3205 (
            .O(N__23978),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    LocalMux I__3204 (
            .O(N__23973),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__3203 (
            .O(N__23968),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__3202 (
            .O(N__23965),
            .I(N__23960));
    InMux I__3201 (
            .O(N__23964),
            .I(N__23955));
    InMux I__3200 (
            .O(N__23963),
            .I(N__23955));
    LocalMux I__3199 (
            .O(N__23960),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    LocalMux I__3198 (
            .O(N__23955),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__3197 (
            .O(N__23950),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__3196 (
            .O(N__23947),
            .I(N__23942));
    InMux I__3195 (
            .O(N__23946),
            .I(N__23937));
    InMux I__3194 (
            .O(N__23945),
            .I(N__23937));
    LocalMux I__3193 (
            .O(N__23942),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    LocalMux I__3192 (
            .O(N__23937),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__3191 (
            .O(N__23932),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__3190 (
            .O(N__23929),
            .I(N__23925));
    CascadeMux I__3189 (
            .O(N__23928),
            .I(N__23921));
    InMux I__3188 (
            .O(N__23925),
            .I(N__23918));
    InMux I__3187 (
            .O(N__23924),
            .I(N__23915));
    InMux I__3186 (
            .O(N__23921),
            .I(N__23912));
    LocalMux I__3185 (
            .O(N__23918),
            .I(N__23909));
    LocalMux I__3184 (
            .O(N__23915),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__3183 (
            .O(N__23912),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__3182 (
            .O(N__23909),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__3181 (
            .O(N__23902),
            .I(bfn_9_23_0_));
    CascadeMux I__3180 (
            .O(N__23899),
            .I(N__23895));
    CascadeMux I__3179 (
            .O(N__23898),
            .I(N__23891));
    InMux I__3178 (
            .O(N__23895),
            .I(N__23888));
    InMux I__3177 (
            .O(N__23894),
            .I(N__23885));
    InMux I__3176 (
            .O(N__23891),
            .I(N__23882));
    LocalMux I__3175 (
            .O(N__23888),
            .I(N__23879));
    LocalMux I__3174 (
            .O(N__23885),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__3173 (
            .O(N__23882),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__3172 (
            .O(N__23879),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__3171 (
            .O(N__23872),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__3170 (
            .O(N__23869),
            .I(N__23865));
    InMux I__3169 (
            .O(N__23868),
            .I(N__23862));
    LocalMux I__3168 (
            .O(N__23865),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    LocalMux I__3167 (
            .O(N__23862),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__3166 (
            .O(N__23857),
            .I(N__23853));
    InMux I__3165 (
            .O(N__23856),
            .I(N__23849));
    InMux I__3164 (
            .O(N__23853),
            .I(N__23846));
    InMux I__3163 (
            .O(N__23852),
            .I(N__23843));
    LocalMux I__3162 (
            .O(N__23849),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__3161 (
            .O(N__23846),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__3160 (
            .O(N__23843),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__3159 (
            .O(N__23836),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__3158 (
            .O(N__23833),
            .I(N__23829));
    InMux I__3157 (
            .O(N__23832),
            .I(N__23825));
    InMux I__3156 (
            .O(N__23829),
            .I(N__23822));
    InMux I__3155 (
            .O(N__23828),
            .I(N__23819));
    LocalMux I__3154 (
            .O(N__23825),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__3153 (
            .O(N__23822),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__3152 (
            .O(N__23819),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__3151 (
            .O(N__23812),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__3150 (
            .O(N__23809),
            .I(N__23804));
    InMux I__3149 (
            .O(N__23808),
            .I(N__23799));
    InMux I__3148 (
            .O(N__23807),
            .I(N__23799));
    LocalMux I__3147 (
            .O(N__23804),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    LocalMux I__3146 (
            .O(N__23799),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__3145 (
            .O(N__23794),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__3144 (
            .O(N__23791),
            .I(N__23787));
    InMux I__3143 (
            .O(N__23790),
            .I(N__23783));
    InMux I__3142 (
            .O(N__23787),
            .I(N__23780));
    InMux I__3141 (
            .O(N__23786),
            .I(N__23777));
    LocalMux I__3140 (
            .O(N__23783),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__3139 (
            .O(N__23780),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__3138 (
            .O(N__23777),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__3137 (
            .O(N__23770),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3136 (
            .O(N__23767),
            .I(N__23762));
    CascadeMux I__3135 (
            .O(N__23766),
            .I(N__23759));
    InMux I__3134 (
            .O(N__23765),
            .I(N__23756));
    InMux I__3133 (
            .O(N__23762),
            .I(N__23751));
    InMux I__3132 (
            .O(N__23759),
            .I(N__23751));
    LocalMux I__3131 (
            .O(N__23756),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    LocalMux I__3130 (
            .O(N__23751),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__3129 (
            .O(N__23746),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__3128 (
            .O(N__23743),
            .I(N__23738));
    InMux I__3127 (
            .O(N__23742),
            .I(N__23733));
    InMux I__3126 (
            .O(N__23741),
            .I(N__23733));
    LocalMux I__3125 (
            .O(N__23738),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    LocalMux I__3124 (
            .O(N__23733),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__3123 (
            .O(N__23728),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__3122 (
            .O(N__23725),
            .I(N__23720));
    InMux I__3121 (
            .O(N__23724),
            .I(N__23715));
    InMux I__3120 (
            .O(N__23723),
            .I(N__23715));
    LocalMux I__3119 (
            .O(N__23720),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    LocalMux I__3118 (
            .O(N__23715),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__3117 (
            .O(N__23710),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3116 (
            .O(N__23707),
            .I(N__23703));
    CascadeMux I__3115 (
            .O(N__23706),
            .I(N__23699));
    InMux I__3114 (
            .O(N__23703),
            .I(N__23696));
    InMux I__3113 (
            .O(N__23702),
            .I(N__23693));
    InMux I__3112 (
            .O(N__23699),
            .I(N__23690));
    LocalMux I__3111 (
            .O(N__23696),
            .I(N__23687));
    LocalMux I__3110 (
            .O(N__23693),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__3109 (
            .O(N__23690),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__3108 (
            .O(N__23687),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__3107 (
            .O(N__23680),
            .I(bfn_9_22_0_));
    CascadeMux I__3106 (
            .O(N__23677),
            .I(N__23673));
    CascadeMux I__3105 (
            .O(N__23676),
            .I(N__23670));
    InMux I__3104 (
            .O(N__23673),
            .I(N__23666));
    InMux I__3103 (
            .O(N__23670),
            .I(N__23663));
    InMux I__3102 (
            .O(N__23669),
            .I(N__23660));
    LocalMux I__3101 (
            .O(N__23666),
            .I(N__23657));
    LocalMux I__3100 (
            .O(N__23663),
            .I(N__23654));
    LocalMux I__3099 (
            .O(N__23660),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__3098 (
            .O(N__23657),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__3097 (
            .O(N__23654),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__3096 (
            .O(N__23647),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__3095 (
            .O(N__23644),
            .I(N__23640));
    InMux I__3094 (
            .O(N__23643),
            .I(N__23636));
    InMux I__3093 (
            .O(N__23640),
            .I(N__23633));
    InMux I__3092 (
            .O(N__23639),
            .I(N__23630));
    LocalMux I__3091 (
            .O(N__23636),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__3090 (
            .O(N__23633),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__3089 (
            .O(N__23630),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__3088 (
            .O(N__23623),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__3087 (
            .O(N__23620),
            .I(N__23615));
    CascadeMux I__3086 (
            .O(N__23619),
            .I(N__23612));
    InMux I__3085 (
            .O(N__23618),
            .I(N__23609));
    InMux I__3084 (
            .O(N__23615),
            .I(N__23604));
    InMux I__3083 (
            .O(N__23612),
            .I(N__23604));
    LocalMux I__3082 (
            .O(N__23609),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    LocalMux I__3081 (
            .O(N__23604),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__3080 (
            .O(N__23599),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__3079 (
            .O(N__23596),
            .I(N__23592));
    CascadeMux I__3078 (
            .O(N__23595),
            .I(N__23589));
    InMux I__3077 (
            .O(N__23592),
            .I(N__23583));
    InMux I__3076 (
            .O(N__23589),
            .I(N__23583));
    InMux I__3075 (
            .O(N__23588),
            .I(N__23580));
    LocalMux I__3074 (
            .O(N__23583),
            .I(N__23577));
    LocalMux I__3073 (
            .O(N__23580),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__3072 (
            .O(N__23577),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__3071 (
            .O(N__23572),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__3070 (
            .O(N__23569),
            .I(N__23565));
    InMux I__3069 (
            .O(N__23568),
            .I(N__23561));
    InMux I__3068 (
            .O(N__23565),
            .I(N__23558));
    InMux I__3067 (
            .O(N__23564),
            .I(N__23555));
    LocalMux I__3066 (
            .O(N__23561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__3065 (
            .O(N__23558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__3064 (
            .O(N__23555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__3063 (
            .O(N__23548),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3062 (
            .O(N__23545),
            .I(N__23541));
    InMux I__3061 (
            .O(N__23544),
            .I(N__23537));
    InMux I__3060 (
            .O(N__23541),
            .I(N__23534));
    InMux I__3059 (
            .O(N__23540),
            .I(N__23531));
    LocalMux I__3058 (
            .O(N__23537),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__3057 (
            .O(N__23534),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__3056 (
            .O(N__23531),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__3055 (
            .O(N__23524),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__3054 (
            .O(N__23521),
            .I(N__23516));
    InMux I__3053 (
            .O(N__23520),
            .I(N__23511));
    InMux I__3052 (
            .O(N__23519),
            .I(N__23511));
    LocalMux I__3051 (
            .O(N__23516),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    LocalMux I__3050 (
            .O(N__23511),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__3049 (
            .O(N__23506),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__3048 (
            .O(N__23503),
            .I(N__23498));
    InMux I__3047 (
            .O(N__23502),
            .I(N__23493));
    InMux I__3046 (
            .O(N__23501),
            .I(N__23493));
    LocalMux I__3045 (
            .O(N__23498),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    LocalMux I__3044 (
            .O(N__23493),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__3043 (
            .O(N__23488),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__3042 (
            .O(N__23485),
            .I(N__23482));
    InMux I__3041 (
            .O(N__23482),
            .I(N__23478));
    CascadeMux I__3040 (
            .O(N__23481),
            .I(N__23474));
    LocalMux I__3039 (
            .O(N__23478),
            .I(N__23471));
    InMux I__3038 (
            .O(N__23477),
            .I(N__23468));
    InMux I__3037 (
            .O(N__23474),
            .I(N__23465));
    Span4Mux_h I__3036 (
            .O(N__23471),
            .I(N__23462));
    LocalMux I__3035 (
            .O(N__23468),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__3034 (
            .O(N__23465),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__3033 (
            .O(N__23462),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__3032 (
            .O(N__23455),
            .I(bfn_9_21_0_));
    CascadeMux I__3031 (
            .O(N__23452),
            .I(N__23448));
    CascadeMux I__3030 (
            .O(N__23451),
            .I(N__23444));
    InMux I__3029 (
            .O(N__23448),
            .I(N__23441));
    InMux I__3028 (
            .O(N__23447),
            .I(N__23438));
    InMux I__3027 (
            .O(N__23444),
            .I(N__23435));
    LocalMux I__3026 (
            .O(N__23441),
            .I(N__23432));
    LocalMux I__3025 (
            .O(N__23438),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__3024 (
            .O(N__23435),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__3023 (
            .O(N__23432),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__3022 (
            .O(N__23425),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__3021 (
            .O(N__23422),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__3020 (
            .O(N__23419),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__3019 (
            .O(N__23416),
            .I(N__23413));
    LocalMux I__3018 (
            .O(N__23413),
            .I(N__23410));
    Span4Mux_h I__3017 (
            .O(N__23410),
            .I(N__23407));
    Odrv4 I__3016 (
            .O(N__23407),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__3015 (
            .O(N__23404),
            .I(N__23401));
    LocalMux I__3014 (
            .O(N__23401),
            .I(\current_shift_inst.control_input_axb_15 ));
    CascadeMux I__3013 (
            .O(N__23398),
            .I(N__23395));
    InMux I__3012 (
            .O(N__23395),
            .I(N__23392));
    LocalMux I__3011 (
            .O(N__23392),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__3010 (
            .O(N__23389),
            .I(N__23386));
    LocalMux I__3009 (
            .O(N__23386),
            .I(N__23383));
    Odrv4 I__3008 (
            .O(N__23383),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__3007 (
            .O(N__23380),
            .I(N__23377));
    LocalMux I__3006 (
            .O(N__23377),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__3005 (
            .O(N__23374),
            .I(N__23371));
    LocalMux I__3004 (
            .O(N__23371),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__3003 (
            .O(N__23368),
            .I(N__23365));
    LocalMux I__3002 (
            .O(N__23365),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__3001 (
            .O(N__23362),
            .I(N__23359));
    LocalMux I__3000 (
            .O(N__23359),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__2999 (
            .O(N__23356),
            .I(N__23353));
    LocalMux I__2998 (
            .O(N__23353),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__2997 (
            .O(N__23350),
            .I(N__23347));
    LocalMux I__2996 (
            .O(N__23347),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__2995 (
            .O(N__23344),
            .I(N__23341));
    LocalMux I__2994 (
            .O(N__23341),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__2993 (
            .O(N__23338),
            .I(N__23335));
    LocalMux I__2992 (
            .O(N__23335),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__2991 (
            .O(N__23332),
            .I(N__23329));
    LocalMux I__2990 (
            .O(N__23329),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__2989 (
            .O(N__23326),
            .I(N__23323));
    LocalMux I__2988 (
            .O(N__23323),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__2987 (
            .O(N__23320),
            .I(N__23317));
    LocalMux I__2986 (
            .O(N__23317),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__2985 (
            .O(N__23314),
            .I(N__23311));
    LocalMux I__2984 (
            .O(N__23311),
            .I(N__23308));
    Span4Mux_v I__2983 (
            .O(N__23308),
            .I(N__23305));
    Odrv4 I__2982 (
            .O(N__23305),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__2981 (
            .O(N__23302),
            .I(N__23299));
    LocalMux I__2980 (
            .O(N__23299),
            .I(N__23296));
    Odrv4 I__2979 (
            .O(N__23296),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__2978 (
            .O(N__23293),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    CascadeMux I__2977 (
            .O(N__23290),
            .I(N__23285));
    InMux I__2976 (
            .O(N__23289),
            .I(N__23282));
    InMux I__2975 (
            .O(N__23288),
            .I(N__23279));
    InMux I__2974 (
            .O(N__23285),
            .I(N__23276));
    LocalMux I__2973 (
            .O(N__23282),
            .I(\current_shift_inst.N_1306_i ));
    LocalMux I__2972 (
            .O(N__23279),
            .I(\current_shift_inst.N_1306_i ));
    LocalMux I__2971 (
            .O(N__23276),
            .I(\current_shift_inst.N_1306_i ));
    InMux I__2970 (
            .O(N__23269),
            .I(N__23266));
    LocalMux I__2969 (
            .O(N__23266),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__2968 (
            .O(N__23263),
            .I(N__23260));
    LocalMux I__2967 (
            .O(N__23260),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__2966 (
            .O(N__23257),
            .I(N__23254));
    LocalMux I__2965 (
            .O(N__23254),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__2964 (
            .O(N__23251),
            .I(N__23248));
    LocalMux I__2963 (
            .O(N__23248),
            .I(\current_shift_inst.control_input_axb_2 ));
    CascadeMux I__2962 (
            .O(N__23245),
            .I(elapsed_time_ns_1_RNI25DN9_0_24_cascade_));
    InMux I__2961 (
            .O(N__23242),
            .I(N__23236));
    InMux I__2960 (
            .O(N__23241),
            .I(N__23236));
    LocalMux I__2959 (
            .O(N__23236),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    InMux I__2958 (
            .O(N__23233),
            .I(N__23228));
    InMux I__2957 (
            .O(N__23232),
            .I(N__23223));
    InMux I__2956 (
            .O(N__23231),
            .I(N__23223));
    LocalMux I__2955 (
            .O(N__23228),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__2954 (
            .O(N__23223),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    CascadeMux I__2953 (
            .O(N__23218),
            .I(N__23214));
    CascadeMux I__2952 (
            .O(N__23217),
            .I(N__23211));
    InMux I__2951 (
            .O(N__23214),
            .I(N__23206));
    InMux I__2950 (
            .O(N__23211),
            .I(N__23206));
    LocalMux I__2949 (
            .O(N__23206),
            .I(N__23203));
    Span4Mux_h I__2948 (
            .O(N__23203),
            .I(N__23200));
    Odrv4 I__2947 (
            .O(N__23200),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__2946 (
            .O(N__23197),
            .I(N__23190));
    InMux I__2945 (
            .O(N__23196),
            .I(N__23190));
    InMux I__2944 (
            .O(N__23195),
            .I(N__23187));
    LocalMux I__2943 (
            .O(N__23190),
            .I(N__23184));
    LocalMux I__2942 (
            .O(N__23187),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__2941 (
            .O(N__23184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    CascadeMux I__2940 (
            .O(N__23179),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ));
    InMux I__2939 (
            .O(N__23176),
            .I(N__23173));
    LocalMux I__2938 (
            .O(N__23173),
            .I(N__23170));
    Span4Mux_v I__2937 (
            .O(N__23170),
            .I(N__23167));
    Odrv4 I__2936 (
            .O(N__23167),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    CascadeMux I__2935 (
            .O(N__23164),
            .I(N__23161));
    InMux I__2934 (
            .O(N__23161),
            .I(N__23158));
    LocalMux I__2933 (
            .O(N__23158),
            .I(N__23155));
    Span4Mux_h I__2932 (
            .O(N__23155),
            .I(N__23152));
    Odrv4 I__2931 (
            .O(N__23152),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    InMux I__2930 (
            .O(N__23149),
            .I(N__23146));
    LocalMux I__2929 (
            .O(N__23146),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__2928 (
            .O(N__23143),
            .I(N__23140));
    LocalMux I__2927 (
            .O(N__23140),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__2926 (
            .O(N__23137),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__2925 (
            .O(N__23134),
            .I(bfn_9_10_0_));
    InMux I__2924 (
            .O(N__23131),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__2923 (
            .O(N__23128),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__2922 (
            .O(N__23125),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__2921 (
            .O(N__23122),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    CascadeMux I__2920 (
            .O(N__23119),
            .I(N__23115));
    InMux I__2919 (
            .O(N__23118),
            .I(N__23112));
    InMux I__2918 (
            .O(N__23115),
            .I(N__23109));
    LocalMux I__2917 (
            .O(N__23112),
            .I(N__23103));
    LocalMux I__2916 (
            .O(N__23109),
            .I(N__23103));
    InMux I__2915 (
            .O(N__23108),
            .I(N__23100));
    Span4Mux_h I__2914 (
            .O(N__23103),
            .I(N__23097));
    LocalMux I__2913 (
            .O(N__23100),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__2912 (
            .O(N__23097),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__2911 (
            .O(N__23092),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__2910 (
            .O(N__23089),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__2909 (
            .O(N__23086),
            .I(N__23082));
    InMux I__2908 (
            .O(N__23085),
            .I(N__23076));
    InMux I__2907 (
            .O(N__23082),
            .I(N__23076));
    InMux I__2906 (
            .O(N__23081),
            .I(N__23073));
    LocalMux I__2905 (
            .O(N__23076),
            .I(N__23070));
    LocalMux I__2904 (
            .O(N__23073),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv12 I__2903 (
            .O(N__23070),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__2902 (
            .O(N__23065),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    CascadeMux I__2901 (
            .O(N__23062),
            .I(N__23057));
    InMux I__2900 (
            .O(N__23061),
            .I(N__23054));
    InMux I__2899 (
            .O(N__23060),
            .I(N__23051));
    InMux I__2898 (
            .O(N__23057),
            .I(N__23048));
    LocalMux I__2897 (
            .O(N__23054),
            .I(N__23045));
    LocalMux I__2896 (
            .O(N__23051),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__2895 (
            .O(N__23048),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__2894 (
            .O(N__23045),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__2893 (
            .O(N__23038),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    CascadeMux I__2892 (
            .O(N__23035),
            .I(N__23032));
    InMux I__2891 (
            .O(N__23032),
            .I(N__23029));
    LocalMux I__2890 (
            .O(N__23029),
            .I(N__23024));
    InMux I__2889 (
            .O(N__23028),
            .I(N__23021));
    InMux I__2888 (
            .O(N__23027),
            .I(N__23018));
    Span4Mux_h I__2887 (
            .O(N__23024),
            .I(N__23015));
    LocalMux I__2886 (
            .O(N__23021),
            .I(N__23012));
    LocalMux I__2885 (
            .O(N__23018),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__2884 (
            .O(N__23015),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__2883 (
            .O(N__23012),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__2882 (
            .O(N__23005),
            .I(bfn_9_9_0_));
    InMux I__2881 (
            .O(N__23002),
            .I(N__22997));
    InMux I__2880 (
            .O(N__23001),
            .I(N__22992));
    InMux I__2879 (
            .O(N__23000),
            .I(N__22992));
    LocalMux I__2878 (
            .O(N__22997),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__2877 (
            .O(N__22992),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__2876 (
            .O(N__22987),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__2875 (
            .O(N__22984),
            .I(N__22979));
    InMux I__2874 (
            .O(N__22983),
            .I(N__22974));
    InMux I__2873 (
            .O(N__22982),
            .I(N__22974));
    LocalMux I__2872 (
            .O(N__22979),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__2871 (
            .O(N__22974),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__2870 (
            .O(N__22969),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__2869 (
            .O(N__22966),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__2868 (
            .O(N__22963),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__2867 (
            .O(N__22960),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__2866 (
            .O(N__22957),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__2865 (
            .O(N__22954),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__2864 (
            .O(N__22951),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__2863 (
            .O(N__22948),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__2862 (
            .O(N__22945),
            .I(bfn_9_8_0_));
    InMux I__2861 (
            .O(N__22942),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__2860 (
            .O(N__22939),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__2859 (
            .O(N__22936),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__2858 (
            .O(N__22933),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__2857 (
            .O(N__22930),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__2856 (
            .O(N__22927),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__2855 (
            .O(N__22924),
            .I(N__22900));
    InMux I__2854 (
            .O(N__22923),
            .I(N__22900));
    InMux I__2853 (
            .O(N__22922),
            .I(N__22900));
    InMux I__2852 (
            .O(N__22921),
            .I(N__22900));
    InMux I__2851 (
            .O(N__22920),
            .I(N__22891));
    InMux I__2850 (
            .O(N__22919),
            .I(N__22891));
    InMux I__2849 (
            .O(N__22918),
            .I(N__22891));
    InMux I__2848 (
            .O(N__22917),
            .I(N__22891));
    InMux I__2847 (
            .O(N__22916),
            .I(N__22868));
    InMux I__2846 (
            .O(N__22915),
            .I(N__22868));
    InMux I__2845 (
            .O(N__22914),
            .I(N__22868));
    InMux I__2844 (
            .O(N__22913),
            .I(N__22868));
    InMux I__2843 (
            .O(N__22912),
            .I(N__22859));
    InMux I__2842 (
            .O(N__22911),
            .I(N__22859));
    InMux I__2841 (
            .O(N__22910),
            .I(N__22859));
    InMux I__2840 (
            .O(N__22909),
            .I(N__22859));
    LocalMux I__2839 (
            .O(N__22900),
            .I(N__22854));
    LocalMux I__2838 (
            .O(N__22891),
            .I(N__22854));
    InMux I__2837 (
            .O(N__22890),
            .I(N__22849));
    InMux I__2836 (
            .O(N__22889),
            .I(N__22849));
    InMux I__2835 (
            .O(N__22888),
            .I(N__22840));
    InMux I__2834 (
            .O(N__22887),
            .I(N__22840));
    InMux I__2833 (
            .O(N__22886),
            .I(N__22840));
    InMux I__2832 (
            .O(N__22885),
            .I(N__22840));
    InMux I__2831 (
            .O(N__22884),
            .I(N__22831));
    InMux I__2830 (
            .O(N__22883),
            .I(N__22831));
    InMux I__2829 (
            .O(N__22882),
            .I(N__22831));
    InMux I__2828 (
            .O(N__22881),
            .I(N__22831));
    InMux I__2827 (
            .O(N__22880),
            .I(N__22822));
    InMux I__2826 (
            .O(N__22879),
            .I(N__22822));
    InMux I__2825 (
            .O(N__22878),
            .I(N__22822));
    InMux I__2824 (
            .O(N__22877),
            .I(N__22822));
    LocalMux I__2823 (
            .O(N__22868),
            .I(N__22817));
    LocalMux I__2822 (
            .O(N__22859),
            .I(N__22817));
    Span4Mux_h I__2821 (
            .O(N__22854),
            .I(N__22814));
    LocalMux I__2820 (
            .O(N__22849),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__2819 (
            .O(N__22840),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__2818 (
            .O(N__22831),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__2817 (
            .O(N__22822),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__2816 (
            .O(N__22817),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__2815 (
            .O(N__22814),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__2814 (
            .O(N__22801),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CEMux I__2813 (
            .O(N__22798),
            .I(N__22794));
    CEMux I__2812 (
            .O(N__22797),
            .I(N__22791));
    LocalMux I__2811 (
            .O(N__22794),
            .I(N__22788));
    LocalMux I__2810 (
            .O(N__22791),
            .I(N__22785));
    Span4Mux_v I__2809 (
            .O(N__22788),
            .I(N__22780));
    Span12Mux_h I__2808 (
            .O(N__22785),
            .I(N__22777));
    CEMux I__2807 (
            .O(N__22784),
            .I(N__22774));
    CEMux I__2806 (
            .O(N__22783),
            .I(N__22771));
    Odrv4 I__2805 (
            .O(N__22780),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    Odrv12 I__2804 (
            .O(N__22777),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    LocalMux I__2803 (
            .O(N__22774),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    LocalMux I__2802 (
            .O(N__22771),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    CascadeMux I__2801 (
            .O(N__22762),
            .I(N__22757));
    InMux I__2800 (
            .O(N__22761),
            .I(N__22753));
    InMux I__2799 (
            .O(N__22760),
            .I(N__22748));
    InMux I__2798 (
            .O(N__22757),
            .I(N__22748));
    InMux I__2797 (
            .O(N__22756),
            .I(N__22745));
    LocalMux I__2796 (
            .O(N__22753),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__2795 (
            .O(N__22748),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__2794 (
            .O(N__22745),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__2793 (
            .O(N__22738),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__2792 (
            .O(N__22735),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__2791 (
            .O(N__22732),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__2790 (
            .O(N__22729),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__2789 (
            .O(N__22726),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__2788 (
            .O(N__22723),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__2787 (
            .O(N__22720),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__2786 (
            .O(N__22717),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__2785 (
            .O(N__22714),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__2784 (
            .O(N__22711),
            .I(bfn_8_24_0_));
    InMux I__2783 (
            .O(N__22708),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__2782 (
            .O(N__22705),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__2781 (
            .O(N__22702),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__2780 (
            .O(N__22699),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__2779 (
            .O(N__22696),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__2778 (
            .O(N__22693),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__2777 (
            .O(N__22690),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__2776 (
            .O(N__22687),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__2775 (
            .O(N__22684),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__2774 (
            .O(N__22681),
            .I(bfn_8_23_0_));
    InMux I__2773 (
            .O(N__22678),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__2772 (
            .O(N__22675),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__2771 (
            .O(N__22672),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__2770 (
            .O(N__22669),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__2769 (
            .O(N__22666),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__2768 (
            .O(N__22663),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__2767 (
            .O(N__22660),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__2766 (
            .O(N__22657),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__2765 (
            .O(N__22654),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__2764 (
            .O(N__22651),
            .I(bfn_8_22_0_));
    InMux I__2763 (
            .O(N__22648),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CEMux I__2762 (
            .O(N__22645),
            .I(N__22639));
    CEMux I__2761 (
            .O(N__22644),
            .I(N__22636));
    CEMux I__2760 (
            .O(N__22643),
            .I(N__22633));
    CEMux I__2759 (
            .O(N__22642),
            .I(N__22630));
    LocalMux I__2758 (
            .O(N__22639),
            .I(N__22624));
    LocalMux I__2757 (
            .O(N__22636),
            .I(N__22624));
    LocalMux I__2756 (
            .O(N__22633),
            .I(N__22621));
    LocalMux I__2755 (
            .O(N__22630),
            .I(N__22618));
    CEMux I__2754 (
            .O(N__22629),
            .I(N__22615));
    Span4Mux_v I__2753 (
            .O(N__22624),
            .I(N__22606));
    Span4Mux_v I__2752 (
            .O(N__22621),
            .I(N__22606));
    Span4Mux_h I__2751 (
            .O(N__22618),
            .I(N__22606));
    LocalMux I__2750 (
            .O(N__22615),
            .I(N__22606));
    Span4Mux_v I__2749 (
            .O(N__22606),
            .I(N__22603));
    Span4Mux_h I__2748 (
            .O(N__22603),
            .I(N__22600));
    Odrv4 I__2747 (
            .O(N__22600),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    CascadeMux I__2746 (
            .O(N__22597),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__2745 (
            .O(N__22594),
            .I(N__22591));
    LocalMux I__2744 (
            .O(N__22591),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__2743 (
            .O(N__22588),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__2742 (
            .O(N__22585),
            .I(bfn_8_21_0_));
    InMux I__2741 (
            .O(N__22582),
            .I(N__22579));
    LocalMux I__2740 (
            .O(N__22579),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__2739 (
            .O(N__22576),
            .I(N__22552));
    InMux I__2738 (
            .O(N__22575),
            .I(N__22552));
    InMux I__2737 (
            .O(N__22574),
            .I(N__22552));
    InMux I__2736 (
            .O(N__22573),
            .I(N__22552));
    InMux I__2735 (
            .O(N__22572),
            .I(N__22533));
    InMux I__2734 (
            .O(N__22571),
            .I(N__22533));
    InMux I__2733 (
            .O(N__22570),
            .I(N__22533));
    InMux I__2732 (
            .O(N__22569),
            .I(N__22533));
    InMux I__2731 (
            .O(N__22568),
            .I(N__22520));
    InMux I__2730 (
            .O(N__22567),
            .I(N__22520));
    InMux I__2729 (
            .O(N__22566),
            .I(N__22520));
    InMux I__2728 (
            .O(N__22565),
            .I(N__22520));
    InMux I__2727 (
            .O(N__22564),
            .I(N__22511));
    InMux I__2726 (
            .O(N__22563),
            .I(N__22511));
    InMux I__2725 (
            .O(N__22562),
            .I(N__22511));
    InMux I__2724 (
            .O(N__22561),
            .I(N__22511));
    LocalMux I__2723 (
            .O(N__22552),
            .I(N__22508));
    InMux I__2722 (
            .O(N__22551),
            .I(N__22499));
    InMux I__2721 (
            .O(N__22550),
            .I(N__22499));
    InMux I__2720 (
            .O(N__22549),
            .I(N__22499));
    InMux I__2719 (
            .O(N__22548),
            .I(N__22499));
    InMux I__2718 (
            .O(N__22547),
            .I(N__22494));
    InMux I__2717 (
            .O(N__22546),
            .I(N__22494));
    InMux I__2716 (
            .O(N__22545),
            .I(N__22485));
    InMux I__2715 (
            .O(N__22544),
            .I(N__22485));
    InMux I__2714 (
            .O(N__22543),
            .I(N__22485));
    InMux I__2713 (
            .O(N__22542),
            .I(N__22485));
    LocalMux I__2712 (
            .O(N__22533),
            .I(N__22482));
    InMux I__2711 (
            .O(N__22532),
            .I(N__22473));
    InMux I__2710 (
            .O(N__22531),
            .I(N__22473));
    InMux I__2709 (
            .O(N__22530),
            .I(N__22473));
    InMux I__2708 (
            .O(N__22529),
            .I(N__22473));
    LocalMux I__2707 (
            .O(N__22520),
            .I(N__22470));
    LocalMux I__2706 (
            .O(N__22511),
            .I(N__22463));
    Span4Mux_h I__2705 (
            .O(N__22508),
            .I(N__22463));
    LocalMux I__2704 (
            .O(N__22499),
            .I(N__22463));
    LocalMux I__2703 (
            .O(N__22494),
            .I(N__22454));
    LocalMux I__2702 (
            .O(N__22485),
            .I(N__22454));
    Span4Mux_v I__2701 (
            .O(N__22482),
            .I(N__22454));
    LocalMux I__2700 (
            .O(N__22473),
            .I(N__22454));
    Span4Mux_v I__2699 (
            .O(N__22470),
            .I(N__22449));
    Span4Mux_v I__2698 (
            .O(N__22463),
            .I(N__22449));
    Span4Mux_v I__2697 (
            .O(N__22454),
            .I(N__22446));
    Odrv4 I__2696 (
            .O(N__22449),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__2695 (
            .O(N__22446),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__2694 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__2693 (
            .O(N__22438),
            .I(N__22435));
    Odrv4 I__2692 (
            .O(N__22435),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__2691 (
            .O(N__22432),
            .I(N__22429));
    LocalMux I__2690 (
            .O(N__22429),
            .I(N__22426));
    Odrv4 I__2689 (
            .O(N__22426),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__2688 (
            .O(N__22423),
            .I(N__22420));
    LocalMux I__2687 (
            .O(N__22420),
            .I(N__22417));
    Span4Mux_v I__2686 (
            .O(N__22417),
            .I(N__22414));
    Odrv4 I__2685 (
            .O(N__22414),
            .I(\current_shift_inst.control_input_axb_7 ));
    CEMux I__2684 (
            .O(N__22411),
            .I(N__22406));
    CEMux I__2683 (
            .O(N__22410),
            .I(N__22403));
    CEMux I__2682 (
            .O(N__22409),
            .I(N__22400));
    LocalMux I__2681 (
            .O(N__22406),
            .I(N__22396));
    LocalMux I__2680 (
            .O(N__22403),
            .I(N__22393));
    LocalMux I__2679 (
            .O(N__22400),
            .I(N__22390));
    CEMux I__2678 (
            .O(N__22399),
            .I(N__22387));
    Span4Mux_v I__2677 (
            .O(N__22396),
            .I(N__22384));
    Span4Mux_v I__2676 (
            .O(N__22393),
            .I(N__22379));
    Span4Mux_h I__2675 (
            .O(N__22390),
            .I(N__22379));
    LocalMux I__2674 (
            .O(N__22387),
            .I(N__22376));
    Span4Mux_v I__2673 (
            .O(N__22384),
            .I(N__22371));
    Span4Mux_v I__2672 (
            .O(N__22379),
            .I(N__22371));
    Span4Mux_v I__2671 (
            .O(N__22376),
            .I(N__22368));
    Odrv4 I__2670 (
            .O(N__22371),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__2669 (
            .O(N__22368),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    InMux I__2668 (
            .O(N__22363),
            .I(N__22357));
    InMux I__2667 (
            .O(N__22362),
            .I(N__22357));
    LocalMux I__2666 (
            .O(N__22357),
            .I(N__22352));
    InMux I__2665 (
            .O(N__22356),
            .I(N__22347));
    InMux I__2664 (
            .O(N__22355),
            .I(N__22347));
    Span12Mux_v I__2663 (
            .O(N__22352),
            .I(N__22344));
    LocalMux I__2662 (
            .O(N__22347),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv12 I__2661 (
            .O(N__22344),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    CascadeMux I__2660 (
            .O(N__22339),
            .I(N__22336));
    InMux I__2659 (
            .O(N__22336),
            .I(N__22326));
    InMux I__2658 (
            .O(N__22335),
            .I(N__22326));
    InMux I__2657 (
            .O(N__22334),
            .I(N__22326));
    InMux I__2656 (
            .O(N__22333),
            .I(N__22323));
    LocalMux I__2655 (
            .O(N__22326),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__2654 (
            .O(N__22323),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__2653 (
            .O(N__22318),
            .I(N__22309));
    InMux I__2652 (
            .O(N__22317),
            .I(N__22309));
    InMux I__2651 (
            .O(N__22316),
            .I(N__22309));
    LocalMux I__2650 (
            .O(N__22309),
            .I(N__22306));
    Span12Mux_v I__2649 (
            .O(N__22306),
            .I(N__22303));
    Odrv12 I__2648 (
            .O(N__22303),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__2647 (
            .O(N__22300),
            .I(N__22297));
    LocalMux I__2646 (
            .O(N__22297),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__2645 (
            .O(N__22294),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__2644 (
            .O(N__22291),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__2643 (
            .O(N__22288),
            .I(N__22285));
    LocalMux I__2642 (
            .O(N__22285),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__2641 (
            .O(N__22282),
            .I(N__22279));
    LocalMux I__2640 (
            .O(N__22279),
            .I(\current_shift_inst.control_input_axb_27 ));
    InMux I__2639 (
            .O(N__22276),
            .I(N__22273));
    LocalMux I__2638 (
            .O(N__22273),
            .I(N__22270));
    Odrv4 I__2637 (
            .O(N__22270),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__2636 (
            .O(N__22267),
            .I(N__22263));
    InMux I__2635 (
            .O(N__22266),
            .I(N__22260));
    LocalMux I__2634 (
            .O(N__22263),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__2633 (
            .O(N__22260),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__2632 (
            .O(N__22255),
            .I(N__22252));
    LocalMux I__2631 (
            .O(N__22252),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__2630 (
            .O(N__22249),
            .I(N__22246));
    LocalMux I__2629 (
            .O(N__22246),
            .I(N__22243));
    Odrv4 I__2628 (
            .O(N__22243),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__2627 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__2626 (
            .O(N__22237),
            .I(N__22234));
    Odrv4 I__2625 (
            .O(N__22234),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__2624 (
            .O(N__22231),
            .I(N__22228));
    LocalMux I__2623 (
            .O(N__22228),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__2622 (
            .O(N__22225),
            .I(N__22222));
    LocalMux I__2621 (
            .O(N__22222),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__2620 (
            .O(N__22219),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__2619 (
            .O(N__22216),
            .I(N__22213));
    LocalMux I__2618 (
            .O(N__22213),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__2617 (
            .O(N__22210),
            .I(\current_shift_inst.control_input_cry_21 ));
    InMux I__2616 (
            .O(N__22207),
            .I(N__22204));
    LocalMux I__2615 (
            .O(N__22204),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__2614 (
            .O(N__22201),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__2613 (
            .O(N__22198),
            .I(N__22195));
    LocalMux I__2612 (
            .O(N__22195),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__2611 (
            .O(N__22192),
            .I(bfn_8_16_0_));
    InMux I__2610 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__2609 (
            .O(N__22186),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__2608 (
            .O(N__22183),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__2607 (
            .O(N__22180),
            .I(N__22177));
    LocalMux I__2606 (
            .O(N__22177),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__2605 (
            .O(N__22174),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__2604 (
            .O(N__22171),
            .I(N__22168));
    LocalMux I__2603 (
            .O(N__22168),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__2602 (
            .O(N__22165),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__2601 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__2600 (
            .O(N__22159),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__2599 (
            .O(N__22156),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__2598 (
            .O(N__22153),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__2597 (
            .O(N__22150),
            .I(N__22147));
    LocalMux I__2596 (
            .O(N__22147),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__2595 (
            .O(N__22144),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__2594 (
            .O(N__22141),
            .I(N__22138));
    LocalMux I__2593 (
            .O(N__22138),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__2592 (
            .O(N__22135),
            .I(\current_shift_inst.control_input_cry_13 ));
    InMux I__2591 (
            .O(N__22132),
            .I(N__22129));
    LocalMux I__2590 (
            .O(N__22129),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__2589 (
            .O(N__22126),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__2588 (
            .O(N__22123),
            .I(N__22120));
    LocalMux I__2587 (
            .O(N__22120),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__2586 (
            .O(N__22117),
            .I(bfn_8_15_0_));
    InMux I__2585 (
            .O(N__22114),
            .I(N__22111));
    LocalMux I__2584 (
            .O(N__22111),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__2583 (
            .O(N__22108),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__2582 (
            .O(N__22105),
            .I(N__22102));
    LocalMux I__2581 (
            .O(N__22102),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__2580 (
            .O(N__22099),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__2579 (
            .O(N__22096),
            .I(N__22093));
    LocalMux I__2578 (
            .O(N__22093),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__2577 (
            .O(N__22090),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__2576 (
            .O(N__22087),
            .I(N__22084));
    LocalMux I__2575 (
            .O(N__22084),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__2574 (
            .O(N__22081),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__2573 (
            .O(N__22078),
            .I(N__22075));
    LocalMux I__2572 (
            .O(N__22075),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__2571 (
            .O(N__22072),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__2570 (
            .O(N__22069),
            .I(N__22066));
    LocalMux I__2569 (
            .O(N__22066),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__2568 (
            .O(N__22063),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__2567 (
            .O(N__22060),
            .I(N__22057));
    LocalMux I__2566 (
            .O(N__22057),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__2565 (
            .O(N__22054),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__2564 (
            .O(N__22051),
            .I(N__22048));
    LocalMux I__2563 (
            .O(N__22048),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__2562 (
            .O(N__22045),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__2561 (
            .O(N__22042),
            .I(N__22039));
    LocalMux I__2560 (
            .O(N__22039),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__2559 (
            .O(N__22036),
            .I(bfn_8_14_0_));
    InMux I__2558 (
            .O(N__22033),
            .I(N__22030));
    LocalMux I__2557 (
            .O(N__22030),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__2556 (
            .O(N__22027),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__2555 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__2554 (
            .O(N__22021),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__2553 (
            .O(N__22018),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__2552 (
            .O(N__22015),
            .I(N__22012));
    LocalMux I__2551 (
            .O(N__22012),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__2550 (
            .O(N__22009),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__2549 (
            .O(N__22006),
            .I(N__22003));
    LocalMux I__2548 (
            .O(N__22003),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    CascadeMux I__2547 (
            .O(N__22000),
            .I(N__21997));
    InMux I__2546 (
            .O(N__21997),
            .I(N__21992));
    InMux I__2545 (
            .O(N__21996),
            .I(N__21989));
    InMux I__2544 (
            .O(N__21995),
            .I(N__21986));
    LocalMux I__2543 (
            .O(N__21992),
            .I(N__21983));
    LocalMux I__2542 (
            .O(N__21989),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__2541 (
            .O(N__21986),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__2540 (
            .O(N__21983),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__2539 (
            .O(N__21976),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__2538 (
            .O(N__21973),
            .I(N__21969));
    InMux I__2537 (
            .O(N__21972),
            .I(N__21966));
    LocalMux I__2536 (
            .O(N__21969),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__2535 (
            .O(N__21966),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__2534 (
            .O(N__21961),
            .I(N__21958));
    InMux I__2533 (
            .O(N__21958),
            .I(N__21953));
    InMux I__2532 (
            .O(N__21957),
            .I(N__21950));
    InMux I__2531 (
            .O(N__21956),
            .I(N__21947));
    LocalMux I__2530 (
            .O(N__21953),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__2529 (
            .O(N__21950),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__2528 (
            .O(N__21947),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__2527 (
            .O(N__21940),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__2526 (
            .O(N__21937),
            .I(N__21933));
    InMux I__2525 (
            .O(N__21936),
            .I(N__21930));
    LocalMux I__2524 (
            .O(N__21933),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__2523 (
            .O(N__21930),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__2522 (
            .O(N__21925),
            .I(N__21920));
    CascadeMux I__2521 (
            .O(N__21924),
            .I(N__21917));
    InMux I__2520 (
            .O(N__21923),
            .I(N__21914));
    InMux I__2519 (
            .O(N__21920),
            .I(N__21909));
    InMux I__2518 (
            .O(N__21917),
            .I(N__21909));
    LocalMux I__2517 (
            .O(N__21914),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__2516 (
            .O(N__21909),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__2515 (
            .O(N__21904),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__2514 (
            .O(N__21901),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__2513 (
            .O(N__21898),
            .I(N__21895));
    LocalMux I__2512 (
            .O(N__21895),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__2511 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__2510 (
            .O(N__21889),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__2509 (
            .O(N__21886),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__2508 (
            .O(N__21883),
            .I(N__21880));
    LocalMux I__2507 (
            .O(N__21880),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__2506 (
            .O(N__21877),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__2505 (
            .O(N__21874),
            .I(N__21871));
    LocalMux I__2504 (
            .O(N__21871),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__2503 (
            .O(N__21868),
            .I(\current_shift_inst.control_input_cry_2 ));
    CascadeMux I__2502 (
            .O(N__21865),
            .I(N__21861));
    CascadeMux I__2501 (
            .O(N__21864),
            .I(N__21858));
    InMux I__2500 (
            .O(N__21861),
            .I(N__21854));
    InMux I__2499 (
            .O(N__21858),
            .I(N__21851));
    InMux I__2498 (
            .O(N__21857),
            .I(N__21848));
    LocalMux I__2497 (
            .O(N__21854),
            .I(N__21845));
    LocalMux I__2496 (
            .O(N__21851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__2495 (
            .O(N__21848),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__2494 (
            .O(N__21845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__2493 (
            .O(N__21838),
            .I(bfn_8_11_0_));
    CascadeMux I__2492 (
            .O(N__21835),
            .I(N__21831));
    CascadeMux I__2491 (
            .O(N__21834),
            .I(N__21828));
    InMux I__2490 (
            .O(N__21831),
            .I(N__21824));
    InMux I__2489 (
            .O(N__21828),
            .I(N__21821));
    InMux I__2488 (
            .O(N__21827),
            .I(N__21818));
    LocalMux I__2487 (
            .O(N__21824),
            .I(N__21815));
    LocalMux I__2486 (
            .O(N__21821),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__2485 (
            .O(N__21818),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__2484 (
            .O(N__21815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__2483 (
            .O(N__21808),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__2482 (
            .O(N__21805),
            .I(N__21802));
    InMux I__2481 (
            .O(N__21802),
            .I(N__21797));
    InMux I__2480 (
            .O(N__21801),
            .I(N__21794));
    InMux I__2479 (
            .O(N__21800),
            .I(N__21791));
    LocalMux I__2478 (
            .O(N__21797),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__2477 (
            .O(N__21794),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__2476 (
            .O(N__21791),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__2475 (
            .O(N__21784),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__2474 (
            .O(N__21781),
            .I(N__21776));
    InMux I__2473 (
            .O(N__21780),
            .I(N__21771));
    InMux I__2472 (
            .O(N__21779),
            .I(N__21771));
    LocalMux I__2471 (
            .O(N__21776),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__2470 (
            .O(N__21771),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__2469 (
            .O(N__21766),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__2468 (
            .O(N__21763),
            .I(N__21760));
    InMux I__2467 (
            .O(N__21760),
            .I(N__21755));
    InMux I__2466 (
            .O(N__21759),
            .I(N__21752));
    InMux I__2465 (
            .O(N__21758),
            .I(N__21749));
    LocalMux I__2464 (
            .O(N__21755),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__2463 (
            .O(N__21752),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__2462 (
            .O(N__21749),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__2461 (
            .O(N__21742),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__2460 (
            .O(N__21739),
            .I(N__21734));
    CascadeMux I__2459 (
            .O(N__21738),
            .I(N__21731));
    InMux I__2458 (
            .O(N__21737),
            .I(N__21728));
    InMux I__2457 (
            .O(N__21734),
            .I(N__21723));
    InMux I__2456 (
            .O(N__21731),
            .I(N__21723));
    LocalMux I__2455 (
            .O(N__21728),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__2454 (
            .O(N__21723),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__2453 (
            .O(N__21718),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__2452 (
            .O(N__21715),
            .I(N__21710));
    InMux I__2451 (
            .O(N__21714),
            .I(N__21705));
    InMux I__2450 (
            .O(N__21713),
            .I(N__21705));
    LocalMux I__2449 (
            .O(N__21710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__2448 (
            .O(N__21705),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__2447 (
            .O(N__21700),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__2446 (
            .O(N__21697),
            .I(N__21692));
    InMux I__2445 (
            .O(N__21696),
            .I(N__21687));
    InMux I__2444 (
            .O(N__21695),
            .I(N__21687));
    LocalMux I__2443 (
            .O(N__21692),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__2442 (
            .O(N__21687),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__2441 (
            .O(N__21682),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__2440 (
            .O(N__21679),
            .I(N__21675));
    CascadeMux I__2439 (
            .O(N__21678),
            .I(N__21672));
    InMux I__2438 (
            .O(N__21675),
            .I(N__21668));
    InMux I__2437 (
            .O(N__21672),
            .I(N__21665));
    InMux I__2436 (
            .O(N__21671),
            .I(N__21662));
    LocalMux I__2435 (
            .O(N__21668),
            .I(N__21659));
    LocalMux I__2434 (
            .O(N__21665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__2433 (
            .O(N__21662),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__2432 (
            .O(N__21659),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__2431 (
            .O(N__21652),
            .I(bfn_8_12_0_));
    CascadeMux I__2430 (
            .O(N__21649),
            .I(N__21645));
    CascadeMux I__2429 (
            .O(N__21648),
            .I(N__21642));
    InMux I__2428 (
            .O(N__21645),
            .I(N__21638));
    InMux I__2427 (
            .O(N__21642),
            .I(N__21635));
    InMux I__2426 (
            .O(N__21641),
            .I(N__21632));
    LocalMux I__2425 (
            .O(N__21638),
            .I(N__21629));
    LocalMux I__2424 (
            .O(N__21635),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__2423 (
            .O(N__21632),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__2422 (
            .O(N__21629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__2421 (
            .O(N__21622),
            .I(bfn_8_10_0_));
    CascadeMux I__2420 (
            .O(N__21619),
            .I(N__21616));
    InMux I__2419 (
            .O(N__21616),
            .I(N__21612));
    CascadeMux I__2418 (
            .O(N__21615),
            .I(N__21609));
    LocalMux I__2417 (
            .O(N__21612),
            .I(N__21605));
    InMux I__2416 (
            .O(N__21609),
            .I(N__21602));
    InMux I__2415 (
            .O(N__21608),
            .I(N__21599));
    Span4Mux_h I__2414 (
            .O(N__21605),
            .I(N__21596));
    LocalMux I__2413 (
            .O(N__21602),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__2412 (
            .O(N__21599),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__2411 (
            .O(N__21596),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__2410 (
            .O(N__21589),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__2409 (
            .O(N__21586),
            .I(N__21583));
    InMux I__2408 (
            .O(N__21583),
            .I(N__21578));
    InMux I__2407 (
            .O(N__21582),
            .I(N__21575));
    InMux I__2406 (
            .O(N__21581),
            .I(N__21572));
    LocalMux I__2405 (
            .O(N__21578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__2404 (
            .O(N__21575),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__2403 (
            .O(N__21572),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__2402 (
            .O(N__21565),
            .I(N__21560));
    CascadeMux I__2401 (
            .O(N__21564),
            .I(N__21556));
    InMux I__2400 (
            .O(N__21563),
            .I(N__21553));
    LocalMux I__2399 (
            .O(N__21560),
            .I(N__21550));
    InMux I__2398 (
            .O(N__21559),
            .I(N__21545));
    InMux I__2397 (
            .O(N__21556),
            .I(N__21545));
    LocalMux I__2396 (
            .O(N__21553),
            .I(N__21542));
    Span4Mux_h I__2395 (
            .O(N__21550),
            .I(N__21539));
    LocalMux I__2394 (
            .O(N__21545),
            .I(N__21536));
    Odrv4 I__2393 (
            .O(N__21542),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__2392 (
            .O(N__21539),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__2391 (
            .O(N__21536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__2390 (
            .O(N__21529),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__2389 (
            .O(N__21526),
            .I(N__21521));
    InMux I__2388 (
            .O(N__21525),
            .I(N__21516));
    InMux I__2387 (
            .O(N__21524),
            .I(N__21516));
    LocalMux I__2386 (
            .O(N__21521),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__2385 (
            .O(N__21516),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__2384 (
            .O(N__21511),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__2383 (
            .O(N__21508),
            .I(N__21505));
    InMux I__2382 (
            .O(N__21505),
            .I(N__21500));
    InMux I__2381 (
            .O(N__21504),
            .I(N__21497));
    InMux I__2380 (
            .O(N__21503),
            .I(N__21494));
    LocalMux I__2379 (
            .O(N__21500),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__2378 (
            .O(N__21497),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__2377 (
            .O(N__21494),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__2376 (
            .O(N__21487),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__2375 (
            .O(N__21484),
            .I(N__21479));
    CascadeMux I__2374 (
            .O(N__21483),
            .I(N__21476));
    InMux I__2373 (
            .O(N__21482),
            .I(N__21473));
    InMux I__2372 (
            .O(N__21479),
            .I(N__21468));
    InMux I__2371 (
            .O(N__21476),
            .I(N__21468));
    LocalMux I__2370 (
            .O(N__21473),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__2369 (
            .O(N__21468),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__2368 (
            .O(N__21463),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__2367 (
            .O(N__21460),
            .I(N__21455));
    InMux I__2366 (
            .O(N__21459),
            .I(N__21450));
    InMux I__2365 (
            .O(N__21458),
            .I(N__21450));
    LocalMux I__2364 (
            .O(N__21455),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__2363 (
            .O(N__21450),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__2362 (
            .O(N__21445),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__2361 (
            .O(N__21442),
            .I(N__21437));
    InMux I__2360 (
            .O(N__21441),
            .I(N__21432));
    InMux I__2359 (
            .O(N__21440),
            .I(N__21432));
    LocalMux I__2358 (
            .O(N__21437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__2357 (
            .O(N__21432),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__2356 (
            .O(N__21427),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__2355 (
            .O(N__21424),
            .I(N__21420));
    InMux I__2354 (
            .O(N__21423),
            .I(N__21416));
    InMux I__2353 (
            .O(N__21420),
            .I(N__21413));
    InMux I__2352 (
            .O(N__21419),
            .I(N__21410));
    LocalMux I__2351 (
            .O(N__21416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__2350 (
            .O(N__21413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__2349 (
            .O(N__21410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__2348 (
            .O(N__21403),
            .I(N__21400));
    InMux I__2347 (
            .O(N__21400),
            .I(N__21396));
    InMux I__2346 (
            .O(N__21399),
            .I(N__21392));
    LocalMux I__2345 (
            .O(N__21396),
            .I(N__21389));
    InMux I__2344 (
            .O(N__21395),
            .I(N__21386));
    LocalMux I__2343 (
            .O(N__21392),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__2342 (
            .O(N__21389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__2341 (
            .O(N__21386),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__2340 (
            .O(N__21379),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__2339 (
            .O(N__21376),
            .I(N__21371));
    InMux I__2338 (
            .O(N__21375),
            .I(N__21366));
    InMux I__2337 (
            .O(N__21374),
            .I(N__21366));
    LocalMux I__2336 (
            .O(N__21371),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__2335 (
            .O(N__21366),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__2334 (
            .O(N__21361),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__2333 (
            .O(N__21358),
            .I(N__21355));
    InMux I__2332 (
            .O(N__21355),
            .I(N__21350));
    InMux I__2331 (
            .O(N__21354),
            .I(N__21347));
    InMux I__2330 (
            .O(N__21353),
            .I(N__21344));
    LocalMux I__2329 (
            .O(N__21350),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__2328 (
            .O(N__21347),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__2327 (
            .O(N__21344),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__2326 (
            .O(N__21337),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__2325 (
            .O(N__21334),
            .I(N__21329));
    CascadeMux I__2324 (
            .O(N__21333),
            .I(N__21326));
    InMux I__2323 (
            .O(N__21332),
            .I(N__21323));
    InMux I__2322 (
            .O(N__21329),
            .I(N__21318));
    InMux I__2321 (
            .O(N__21326),
            .I(N__21318));
    LocalMux I__2320 (
            .O(N__21323),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__2319 (
            .O(N__21318),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__2318 (
            .O(N__21313),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__2317 (
            .O(N__21310),
            .I(N__21307));
    InMux I__2316 (
            .O(N__21307),
            .I(N__21302));
    InMux I__2315 (
            .O(N__21306),
            .I(N__21299));
    InMux I__2314 (
            .O(N__21305),
            .I(N__21296));
    LocalMux I__2313 (
            .O(N__21302),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__2312 (
            .O(N__21299),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__2311 (
            .O(N__21296),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__2310 (
            .O(N__21289),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__2309 (
            .O(N__21286),
            .I(N__21281));
    InMux I__2308 (
            .O(N__21285),
            .I(N__21276));
    InMux I__2307 (
            .O(N__21284),
            .I(N__21276));
    LocalMux I__2306 (
            .O(N__21281),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__2305 (
            .O(N__21276),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__2304 (
            .O(N__21271),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__2303 (
            .O(N__21268),
            .I(N__21263));
    InMux I__2302 (
            .O(N__21267),
            .I(N__21258));
    InMux I__2301 (
            .O(N__21266),
            .I(N__21258));
    LocalMux I__2300 (
            .O(N__21263),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__2299 (
            .O(N__21258),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__2298 (
            .O(N__21253),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__2297 (
            .O(N__21250),
            .I(N__21246));
    InMux I__2296 (
            .O(N__21249),
            .I(N__21243));
    LocalMux I__2295 (
            .O(N__21246),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    LocalMux I__2294 (
            .O(N__21243),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__2293 (
            .O(N__21238),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    InMux I__2292 (
            .O(N__21235),
            .I(N__21231));
    InMux I__2291 (
            .O(N__21234),
            .I(N__21228));
    LocalMux I__2290 (
            .O(N__21231),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    LocalMux I__2289 (
            .O(N__21228),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__2288 (
            .O(N__21223),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__2287 (
            .O(N__21220),
            .I(N__21214));
    InMux I__2286 (
            .O(N__21219),
            .I(N__21214));
    LocalMux I__2285 (
            .O(N__21214),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__2284 (
            .O(N__21211),
            .I(N__21207));
    CascadeMux I__2283 (
            .O(N__21210),
            .I(N__21204));
    InMux I__2282 (
            .O(N__21207),
            .I(N__21199));
    InMux I__2281 (
            .O(N__21204),
            .I(N__21199));
    LocalMux I__2280 (
            .O(N__21199),
            .I(N__21196));
    Odrv4 I__2279 (
            .O(N__21196),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__2278 (
            .O(N__21193),
            .I(N__21190));
    LocalMux I__2277 (
            .O(N__21190),
            .I(N__21187));
    Span4Mux_s3_h I__2276 (
            .O(N__21187),
            .I(N__21183));
    InMux I__2275 (
            .O(N__21186),
            .I(N__21180));
    Span4Mux_h I__2274 (
            .O(N__21183),
            .I(N__21177));
    LocalMux I__2273 (
            .O(N__21180),
            .I(N__21174));
    Sp12to4 I__2272 (
            .O(N__21177),
            .I(N__21171));
    Odrv12 I__2271 (
            .O(N__21174),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv12 I__2270 (
            .O(N__21171),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__2269 (
            .O(N__21166),
            .I(N__21158));
    InMux I__2268 (
            .O(N__21165),
            .I(N__21158));
    InMux I__2267 (
            .O(N__21164),
            .I(N__21155));
    InMux I__2266 (
            .O(N__21163),
            .I(N__21152));
    LocalMux I__2265 (
            .O(N__21158),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__2264 (
            .O(N__21155),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__2263 (
            .O(N__21152),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__2262 (
            .O(N__21145),
            .I(N__21139));
    InMux I__2261 (
            .O(N__21144),
            .I(N__21134));
    InMux I__2260 (
            .O(N__21143),
            .I(N__21134));
    InMux I__2259 (
            .O(N__21142),
            .I(N__21131));
    LocalMux I__2258 (
            .O(N__21139),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__2257 (
            .O(N__21134),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__2256 (
            .O(N__21131),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    IoInMux I__2255 (
            .O(N__21124),
            .I(N__21121));
    LocalMux I__2254 (
            .O(N__21121),
            .I(N__21118));
    Span4Mux_s0_v I__2253 (
            .O(N__21118),
            .I(N__21115));
    Span4Mux_h I__2252 (
            .O(N__21115),
            .I(N__21112));
    Span4Mux_v I__2251 (
            .O(N__21112),
            .I(N__21109));
    Odrv4 I__2250 (
            .O(N__21109),
            .I(\current_shift_inst.timer_s1.N_161_i ));
    ClkMux I__2249 (
            .O(N__21106),
            .I(N__21103));
    GlobalMux I__2248 (
            .O(N__21103),
            .I(N__21100));
    gio2CtrlBuf I__2247 (
            .O(N__21100),
            .I(delay_hc_input_c_g));
    InMux I__2246 (
            .O(N__21097),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__2245 (
            .O(N__21094),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__2244 (
            .O(N__21091),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__2243 (
            .O(N__21088),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__2242 (
            .O(N__21085),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__2241 (
            .O(N__21082),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__2240 (
            .O(N__21079),
            .I(N__21076));
    LocalMux I__2239 (
            .O(N__21076),
            .I(N__21073));
    Span4Mux_s3_h I__2238 (
            .O(N__21073),
            .I(N__21070));
    Span4Mux_v I__2237 (
            .O(N__21070),
            .I(N__21067));
    Span4Mux_v I__2236 (
            .O(N__21067),
            .I(N__21063));
    InMux I__2235 (
            .O(N__21066),
            .I(N__21060));
    Span4Mux_h I__2234 (
            .O(N__21063),
            .I(N__21057));
    LocalMux I__2233 (
            .O(N__21060),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv4 I__2232 (
            .O(N__21057),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__2231 (
            .O(N__21052),
            .I(N__21049));
    LocalMux I__2230 (
            .O(N__21049),
            .I(N__21045));
    InMux I__2229 (
            .O(N__21048),
            .I(N__21042));
    Span12Mux_v I__2228 (
            .O(N__21045),
            .I(N__21039));
    LocalMux I__2227 (
            .O(N__21042),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    Odrv12 I__2226 (
            .O(N__21039),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__2225 (
            .O(N__21034),
            .I(N__21031));
    LocalMux I__2224 (
            .O(N__21031),
            .I(N__21027));
    InMux I__2223 (
            .O(N__21030),
            .I(N__21024));
    Span4Mux_h I__2222 (
            .O(N__21027),
            .I(N__21021));
    LocalMux I__2221 (
            .O(N__21024),
            .I(N__21018));
    Span4Mux_v I__2220 (
            .O(N__21021),
            .I(N__21015));
    Span4Mux_v I__2219 (
            .O(N__21018),
            .I(N__21010));
    Span4Mux_v I__2218 (
            .O(N__21015),
            .I(N__21010));
    Odrv4 I__2217 (
            .O(N__21010),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__2216 (
            .O(N__21007),
            .I(N__21003));
    InMux I__2215 (
            .O(N__21006),
            .I(N__21000));
    LocalMux I__2214 (
            .O(N__21003),
            .I(N__20997));
    LocalMux I__2213 (
            .O(N__21000),
            .I(N__20994));
    Span12Mux_s7_h I__2212 (
            .O(N__20997),
            .I(N__20991));
    Odrv4 I__2211 (
            .O(N__20994),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv12 I__2210 (
            .O(N__20991),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__2209 (
            .O(N__20986),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__2208 (
            .O(N__20983),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__2207 (
            .O(N__20980),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__2206 (
            .O(N__20977),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__2205 (
            .O(N__20974),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__2204 (
            .O(N__20971),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__2203 (
            .O(N__20968),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__2202 (
            .O(N__20965),
            .I(bfn_7_17_0_));
    InMux I__2201 (
            .O(N__20962),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__2200 (
            .O(N__20959),
            .I(bfn_7_15_0_));
    InMux I__2199 (
            .O(N__20956),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__2198 (
            .O(N__20953),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__2197 (
            .O(N__20950),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__2196 (
            .O(N__20947),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__2195 (
            .O(N__20944),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__2194 (
            .O(N__20941),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__2193 (
            .O(N__20938),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__2192 (
            .O(N__20935),
            .I(bfn_7_16_0_));
    InMux I__2191 (
            .O(N__20932),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__2190 (
            .O(N__20929),
            .I(N__20926));
    LocalMux I__2189 (
            .O(N__20926),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__2188 (
            .O(N__20923),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__2187 (
            .O(N__20920),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__2186 (
            .O(N__20917),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__2185 (
            .O(N__20914),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__2184 (
            .O(N__20911),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__2183 (
            .O(N__20908),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__2182 (
            .O(N__20905),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__2181 (
            .O(N__20902),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__2180 (
            .O(N__20899),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__2179 (
            .O(N__20896),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__2178 (
            .O(N__20893),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__2177 (
            .O(N__20890),
            .I(bfn_7_13_0_));
    InMux I__2176 (
            .O(N__20887),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__2175 (
            .O(N__20884),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__2174 (
            .O(N__20881),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__2173 (
            .O(N__20878),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__2172 (
            .O(N__20875),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__2171 (
            .O(N__20872),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__2170 (
            .O(N__20869),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__2169 (
            .O(N__20866),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__2168 (
            .O(N__20863),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__2167 (
            .O(N__20860),
            .I(bfn_7_12_0_));
    InMux I__2166 (
            .O(N__20857),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__2165 (
            .O(N__20854),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__2164 (
            .O(N__20851),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__2163 (
            .O(N__20848),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__2162 (
            .O(N__20845),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__2161 (
            .O(N__20842),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__2160 (
            .O(N__20839),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__2159 (
            .O(N__20836),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__2158 (
            .O(N__20833),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__2157 (
            .O(N__20830),
            .I(bfn_7_11_0_));
    InMux I__2156 (
            .O(N__20827),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__2155 (
            .O(N__20824),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__2154 (
            .O(N__20821),
            .I(N__20818));
    LocalMux I__2153 (
            .O(N__20818),
            .I(N__20814));
    InMux I__2152 (
            .O(N__20817),
            .I(N__20810));
    Span4Mux_h I__2151 (
            .O(N__20814),
            .I(N__20807));
    InMux I__2150 (
            .O(N__20813),
            .I(N__20804));
    LocalMux I__2149 (
            .O(N__20810),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__2148 (
            .O(N__20807),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__2147 (
            .O(N__20804),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    CascadeMux I__2146 (
            .O(N__20797),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__2145 (
            .O(N__20794),
            .I(N__20791));
    LocalMux I__2144 (
            .O(N__20791),
            .I(N__20788));
    Odrv12 I__2143 (
            .O(N__20788),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__2142 (
            .O(N__20785),
            .I(bfn_7_10_0_));
    InMux I__2141 (
            .O(N__20782),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__2140 (
            .O(N__20779),
            .I(N__20773));
    InMux I__2139 (
            .O(N__20778),
            .I(N__20773));
    LocalMux I__2138 (
            .O(N__20773),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__2137 (
            .O(N__20770),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    InMux I__2136 (
            .O(N__20767),
            .I(N__20764));
    LocalMux I__2135 (
            .O(N__20764),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__2134 (
            .O(N__20761),
            .I(N__20758));
    LocalMux I__2133 (
            .O(N__20758),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    CascadeMux I__2132 (
            .O(N__20755),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__2131 (
            .O(N__20752),
            .I(N__20748));
    InMux I__2130 (
            .O(N__20751),
            .I(N__20745));
    LocalMux I__2129 (
            .O(N__20748),
            .I(N__20740));
    LocalMux I__2128 (
            .O(N__20745),
            .I(N__20740));
    Odrv4 I__2127 (
            .O(N__20740),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__2126 (
            .O(N__20737),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__2125 (
            .O(N__20734),
            .I(N__20731));
    LocalMux I__2124 (
            .O(N__20731),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__2123 (
            .O(N__20728),
            .I(N__20725));
    LocalMux I__2122 (
            .O(N__20725),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    CascadeMux I__2121 (
            .O(N__20722),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    CascadeMux I__2120 (
            .O(N__20719),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    InMux I__2119 (
            .O(N__20716),
            .I(N__20713));
    LocalMux I__2118 (
            .O(N__20713),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__2117 (
            .O(N__20710),
            .I(N__20707));
    LocalMux I__2116 (
            .O(N__20707),
            .I(N__20704));
    Odrv12 I__2115 (
            .O(N__20704),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2114 (
            .O(N__20701),
            .I(N__20698));
    LocalMux I__2113 (
            .O(N__20698),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__2112 (
            .O(N__20695),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    CascadeMux I__2111 (
            .O(N__20692),
            .I(N__20682));
    CascadeMux I__2110 (
            .O(N__20691),
            .I(N__20679));
    CascadeMux I__2109 (
            .O(N__20690),
            .I(N__20667));
    CascadeMux I__2108 (
            .O(N__20689),
            .I(N__20664));
    CascadeMux I__2107 (
            .O(N__20688),
            .I(N__20661));
    CascadeMux I__2106 (
            .O(N__20687),
            .I(N__20657));
    InMux I__2105 (
            .O(N__20686),
            .I(N__20638));
    InMux I__2104 (
            .O(N__20685),
            .I(N__20638));
    InMux I__2103 (
            .O(N__20682),
            .I(N__20638));
    InMux I__2102 (
            .O(N__20679),
            .I(N__20638));
    InMux I__2101 (
            .O(N__20678),
            .I(N__20638));
    InMux I__2100 (
            .O(N__20677),
            .I(N__20633));
    InMux I__2099 (
            .O(N__20676),
            .I(N__20633));
    InMux I__2098 (
            .O(N__20675),
            .I(N__20624));
    InMux I__2097 (
            .O(N__20674),
            .I(N__20624));
    InMux I__2096 (
            .O(N__20673),
            .I(N__20624));
    InMux I__2095 (
            .O(N__20672),
            .I(N__20624));
    CascadeMux I__2094 (
            .O(N__20671),
            .I(N__20620));
    CascadeMux I__2093 (
            .O(N__20670),
            .I(N__20617));
    InMux I__2092 (
            .O(N__20667),
            .I(N__20606));
    InMux I__2091 (
            .O(N__20664),
            .I(N__20606));
    InMux I__2090 (
            .O(N__20661),
            .I(N__20606));
    InMux I__2089 (
            .O(N__20660),
            .I(N__20606));
    InMux I__2088 (
            .O(N__20657),
            .I(N__20599));
    InMux I__2087 (
            .O(N__20656),
            .I(N__20599));
    InMux I__2086 (
            .O(N__20655),
            .I(N__20599));
    InMux I__2085 (
            .O(N__20654),
            .I(N__20594));
    InMux I__2084 (
            .O(N__20653),
            .I(N__20583));
    InMux I__2083 (
            .O(N__20652),
            .I(N__20583));
    InMux I__2082 (
            .O(N__20651),
            .I(N__20583));
    InMux I__2081 (
            .O(N__20650),
            .I(N__20583));
    InMux I__2080 (
            .O(N__20649),
            .I(N__20583));
    LocalMux I__2079 (
            .O(N__20638),
            .I(N__20580));
    LocalMux I__2078 (
            .O(N__20633),
            .I(N__20575));
    LocalMux I__2077 (
            .O(N__20624),
            .I(N__20575));
    InMux I__2076 (
            .O(N__20623),
            .I(N__20572));
    InMux I__2075 (
            .O(N__20620),
            .I(N__20563));
    InMux I__2074 (
            .O(N__20617),
            .I(N__20563));
    InMux I__2073 (
            .O(N__20616),
            .I(N__20563));
    InMux I__2072 (
            .O(N__20615),
            .I(N__20563));
    LocalMux I__2071 (
            .O(N__20606),
            .I(N__20558));
    LocalMux I__2070 (
            .O(N__20599),
            .I(N__20558));
    InMux I__2069 (
            .O(N__20598),
            .I(N__20555));
    InMux I__2068 (
            .O(N__20597),
            .I(N__20552));
    LocalMux I__2067 (
            .O(N__20594),
            .I(N__20547));
    LocalMux I__2066 (
            .O(N__20583),
            .I(N__20547));
    Span4Mux_v I__2065 (
            .O(N__20580),
            .I(N__20542));
    Span4Mux_h I__2064 (
            .O(N__20575),
            .I(N__20542));
    LocalMux I__2063 (
            .O(N__20572),
            .I(N__20535));
    LocalMux I__2062 (
            .O(N__20563),
            .I(N__20535));
    Sp12to4 I__2061 (
            .O(N__20558),
            .I(N__20535));
    LocalMux I__2060 (
            .O(N__20555),
            .I(N__20528));
    LocalMux I__2059 (
            .O(N__20552),
            .I(N__20528));
    Span4Mux_h I__2058 (
            .O(N__20547),
            .I(N__20528));
    Odrv4 I__2057 (
            .O(N__20542),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv12 I__2056 (
            .O(N__20535),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2055 (
            .O(N__20528),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    InMux I__2054 (
            .O(N__20521),
            .I(N__20518));
    LocalMux I__2053 (
            .O(N__20518),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    CascadeMux I__2052 (
            .O(N__20515),
            .I(N__20512));
    InMux I__2051 (
            .O(N__20512),
            .I(N__20509));
    LocalMux I__2050 (
            .O(N__20509),
            .I(N__20506));
    Odrv4 I__2049 (
            .O(N__20506),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2048 (
            .O(N__20503),
            .I(N__20500));
    LocalMux I__2047 (
            .O(N__20500),
            .I(N__20497));
    Odrv4 I__2046 (
            .O(N__20497),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__2045 (
            .O(N__20494),
            .I(N__20491));
    InMux I__2044 (
            .O(N__20491),
            .I(N__20488));
    LocalMux I__2043 (
            .O(N__20488),
            .I(N__20485));
    Span4Mux_h I__2042 (
            .O(N__20485),
            .I(N__20482));
    Odrv4 I__2041 (
            .O(N__20482),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__2040 (
            .O(N__20479),
            .I(N__20476));
    InMux I__2039 (
            .O(N__20476),
            .I(N__20473));
    LocalMux I__2038 (
            .O(N__20473),
            .I(N__20470));
    Span4Mux_h I__2037 (
            .O(N__20470),
            .I(N__20467));
    Odrv4 I__2036 (
            .O(N__20467),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__2035 (
            .O(N__20464),
            .I(N__20461));
    LocalMux I__2034 (
            .O(N__20461),
            .I(N__20458));
    Span4Mux_h I__2033 (
            .O(N__20458),
            .I(N__20455));
    Odrv4 I__2032 (
            .O(N__20455),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__2031 (
            .O(N__20452),
            .I(N__20449));
    InMux I__2030 (
            .O(N__20449),
            .I(N__20446));
    LocalMux I__2029 (
            .O(N__20446),
            .I(N__20443));
    Span4Mux_h I__2028 (
            .O(N__20443),
            .I(N__20440));
    Odrv4 I__2027 (
            .O(N__20440),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__2026 (
            .O(N__20437),
            .I(N__20414));
    CascadeMux I__2025 (
            .O(N__20436),
            .I(N__20411));
    CascadeMux I__2024 (
            .O(N__20435),
            .I(N__20408));
    CascadeMux I__2023 (
            .O(N__20434),
            .I(N__20405));
    InMux I__2022 (
            .O(N__20433),
            .I(N__20395));
    InMux I__2021 (
            .O(N__20432),
            .I(N__20386));
    InMux I__2020 (
            .O(N__20431),
            .I(N__20386));
    InMux I__2019 (
            .O(N__20430),
            .I(N__20386));
    InMux I__2018 (
            .O(N__20429),
            .I(N__20386));
    CascadeMux I__2017 (
            .O(N__20428),
            .I(N__20382));
    CascadeMux I__2016 (
            .O(N__20427),
            .I(N__20379));
    CascadeMux I__2015 (
            .O(N__20426),
            .I(N__20374));
    CascadeMux I__2014 (
            .O(N__20425),
            .I(N__20371));
    InMux I__2013 (
            .O(N__20424),
            .I(N__20364));
    InMux I__2012 (
            .O(N__20423),
            .I(N__20364));
    InMux I__2011 (
            .O(N__20422),
            .I(N__20364));
    InMux I__2010 (
            .O(N__20421),
            .I(N__20355));
    InMux I__2009 (
            .O(N__20420),
            .I(N__20355));
    InMux I__2008 (
            .O(N__20419),
            .I(N__20355));
    InMux I__2007 (
            .O(N__20418),
            .I(N__20355));
    InMux I__2006 (
            .O(N__20417),
            .I(N__20352));
    InMux I__2005 (
            .O(N__20414),
            .I(N__20349));
    InMux I__2004 (
            .O(N__20411),
            .I(N__20338));
    InMux I__2003 (
            .O(N__20408),
            .I(N__20338));
    InMux I__2002 (
            .O(N__20405),
            .I(N__20338));
    InMux I__2001 (
            .O(N__20404),
            .I(N__20338));
    InMux I__2000 (
            .O(N__20403),
            .I(N__20338));
    InMux I__1999 (
            .O(N__20402),
            .I(N__20327));
    InMux I__1998 (
            .O(N__20401),
            .I(N__20327));
    InMux I__1997 (
            .O(N__20400),
            .I(N__20327));
    InMux I__1996 (
            .O(N__20399),
            .I(N__20327));
    InMux I__1995 (
            .O(N__20398),
            .I(N__20327));
    LocalMux I__1994 (
            .O(N__20395),
            .I(N__20324));
    LocalMux I__1993 (
            .O(N__20386),
            .I(N__20321));
    InMux I__1992 (
            .O(N__20385),
            .I(N__20318));
    InMux I__1991 (
            .O(N__20382),
            .I(N__20313));
    InMux I__1990 (
            .O(N__20379),
            .I(N__20313));
    InMux I__1989 (
            .O(N__20378),
            .I(N__20304));
    InMux I__1988 (
            .O(N__20377),
            .I(N__20304));
    InMux I__1987 (
            .O(N__20374),
            .I(N__20304));
    InMux I__1986 (
            .O(N__20371),
            .I(N__20304));
    LocalMux I__1985 (
            .O(N__20364),
            .I(N__20299));
    LocalMux I__1984 (
            .O(N__20355),
            .I(N__20299));
    LocalMux I__1983 (
            .O(N__20352),
            .I(N__20286));
    LocalMux I__1982 (
            .O(N__20349),
            .I(N__20286));
    LocalMux I__1981 (
            .O(N__20338),
            .I(N__20286));
    LocalMux I__1980 (
            .O(N__20327),
            .I(N__20286));
    Span4Mux_v I__1979 (
            .O(N__20324),
            .I(N__20286));
    Span4Mux_h I__1978 (
            .O(N__20321),
            .I(N__20286));
    LocalMux I__1977 (
            .O(N__20318),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__1976 (
            .O(N__20313),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__1975 (
            .O(N__20304),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv12 I__1974 (
            .O(N__20299),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__1973 (
            .O(N__20286),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    InMux I__1972 (
            .O(N__20275),
            .I(N__20272));
    LocalMux I__1971 (
            .O(N__20272),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    CascadeMux I__1970 (
            .O(N__20269),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__1969 (
            .O(N__20266),
            .I(N__20263));
    LocalMux I__1968 (
            .O(N__20263),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__1967 (
            .O(N__20260),
            .I(N__20257));
    LocalMux I__1966 (
            .O(N__20257),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    CascadeMux I__1965 (
            .O(N__20254),
            .I(N__20251));
    InMux I__1964 (
            .O(N__20251),
            .I(N__20248));
    LocalMux I__1963 (
            .O(N__20248),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    CascadeMux I__1962 (
            .O(N__20245),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    InMux I__1961 (
            .O(N__20242),
            .I(N__20239));
    LocalMux I__1960 (
            .O(N__20239),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__1959 (
            .O(N__20236),
            .I(N__20232));
    CascadeMux I__1958 (
            .O(N__20235),
            .I(N__20229));
    InMux I__1957 (
            .O(N__20232),
            .I(N__20226));
    InMux I__1956 (
            .O(N__20229),
            .I(N__20223));
    LocalMux I__1955 (
            .O(N__20226),
            .I(N__20218));
    LocalMux I__1954 (
            .O(N__20223),
            .I(N__20218));
    Span4Mux_h I__1953 (
            .O(N__20218),
            .I(N__20215));
    Odrv4 I__1952 (
            .O(N__20215),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    InMux I__1951 (
            .O(N__20212),
            .I(N__20209));
    LocalMux I__1950 (
            .O(N__20209),
            .I(N__20206));
    Odrv4 I__1949 (
            .O(N__20206),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    CascadeMux I__1948 (
            .O(N__20203),
            .I(N__20200));
    InMux I__1947 (
            .O(N__20200),
            .I(N__20197));
    LocalMux I__1946 (
            .O(N__20197),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__1945 (
            .O(N__20194),
            .I(N__20191));
    LocalMux I__1944 (
            .O(N__20191),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__1943 (
            .O(N__20188),
            .I(N__20185));
    LocalMux I__1942 (
            .O(N__20185),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__1941 (
            .O(N__20182),
            .I(N__20179));
    LocalMux I__1940 (
            .O(N__20179),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__1939 (
            .O(N__20176),
            .I(N__20173));
    InMux I__1938 (
            .O(N__20173),
            .I(N__20170));
    LocalMux I__1937 (
            .O(N__20170),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__1936 (
            .O(N__20167),
            .I(N__20164));
    LocalMux I__1935 (
            .O(N__20164),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__1934 (
            .O(N__20161),
            .I(N__20158));
    InMux I__1933 (
            .O(N__20158),
            .I(N__20155));
    LocalMux I__1932 (
            .O(N__20155),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    CascadeMux I__1931 (
            .O(N__20152),
            .I(N__20149));
    InMux I__1930 (
            .O(N__20149),
            .I(N__20146));
    LocalMux I__1929 (
            .O(N__20146),
            .I(N__20143));
    Odrv4 I__1928 (
            .O(N__20143),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__1927 (
            .O(N__20140),
            .I(N__20137));
    LocalMux I__1926 (
            .O(N__20137),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__1925 (
            .O(N__20134),
            .I(N__20131));
    LocalMux I__1924 (
            .O(N__20131),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__1923 (
            .O(N__20128),
            .I(N__20125));
    LocalMux I__1922 (
            .O(N__20125),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    CascadeMux I__1921 (
            .O(N__20122),
            .I(N__20119));
    InMux I__1920 (
            .O(N__20119),
            .I(N__20116));
    LocalMux I__1919 (
            .O(N__20116),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__1918 (
            .O(N__20113),
            .I(N__20110));
    LocalMux I__1917 (
            .O(N__20110),
            .I(N__20107));
    Odrv4 I__1916 (
            .O(N__20107),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__1915 (
            .O(N__20104),
            .I(N__20101));
    LocalMux I__1914 (
            .O(N__20101),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    CascadeMux I__1913 (
            .O(N__20098),
            .I(N__20095));
    InMux I__1912 (
            .O(N__20095),
            .I(N__20092));
    LocalMux I__1911 (
            .O(N__20092),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__1910 (
            .O(N__20089),
            .I(N__20086));
    LocalMux I__1909 (
            .O(N__20086),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__1908 (
            .O(N__20083),
            .I(N__20080));
    InMux I__1907 (
            .O(N__20080),
            .I(N__20077));
    LocalMux I__1906 (
            .O(N__20077),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__1905 (
            .O(N__20074),
            .I(N__20071));
    LocalMux I__1904 (
            .O(N__20071),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    CascadeMux I__1903 (
            .O(N__20068),
            .I(N__20065));
    InMux I__1902 (
            .O(N__20065),
            .I(N__20062));
    LocalMux I__1901 (
            .O(N__20062),
            .I(N__20059));
    Span4Mux_v I__1900 (
            .O(N__20059),
            .I(N__20056));
    Odrv4 I__1899 (
            .O(N__20056),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1898 (
            .O(N__20053),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__1897 (
            .O(N__20050),
            .I(N__20047));
    InMux I__1896 (
            .O(N__20047),
            .I(N__20044));
    LocalMux I__1895 (
            .O(N__20044),
            .I(N__20041));
    Odrv4 I__1894 (
            .O(N__20041),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1893 (
            .O(N__20038),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__1892 (
            .O(N__20035),
            .I(N__20032));
    InMux I__1891 (
            .O(N__20032),
            .I(N__20029));
    LocalMux I__1890 (
            .O(N__20029),
            .I(N__20026));
    Span4Mux_v I__1889 (
            .O(N__20026),
            .I(N__20023));
    Odrv4 I__1888 (
            .O(N__20023),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1887 (
            .O(N__20020),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__1886 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__1885 (
            .O(N__20014),
            .I(N__20011));
    Odrv4 I__1884 (
            .O(N__20011),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__1883 (
            .O(N__20008),
            .I(N__20005));
    InMux I__1882 (
            .O(N__20005),
            .I(N__20002));
    LocalMux I__1881 (
            .O(N__20002),
            .I(N__19999));
    Span4Mux_v I__1880 (
            .O(N__19999),
            .I(N__19996));
    Odrv4 I__1879 (
            .O(N__19996),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__1878 (
            .O(N__19993),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    CascadeMux I__1877 (
            .O(N__19990),
            .I(N__19987));
    InMux I__1876 (
            .O(N__19987),
            .I(N__19984));
    LocalMux I__1875 (
            .O(N__19984),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__1874 (
            .O(N__19981),
            .I(N__19978));
    LocalMux I__1873 (
            .O(N__19978),
            .I(N__19975));
    Odrv12 I__1872 (
            .O(N__19975),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__1871 (
            .O(N__19972),
            .I(N__19969));
    LocalMux I__1870 (
            .O(N__19969),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__1869 (
            .O(N__19966),
            .I(N__19963));
    InMux I__1868 (
            .O(N__19963),
            .I(N__19960));
    LocalMux I__1867 (
            .O(N__19960),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__1866 (
            .O(N__19957),
            .I(N__19954));
    LocalMux I__1865 (
            .O(N__19954),
            .I(N__19951));
    Odrv4 I__1864 (
            .O(N__19951),
            .I(N_39_i_i));
    CascadeMux I__1863 (
            .O(N__19948),
            .I(N__19945));
    InMux I__1862 (
            .O(N__19945),
            .I(N__19942));
    LocalMux I__1861 (
            .O(N__19942),
            .I(N__19939));
    Odrv4 I__1860 (
            .O(N__19939),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1859 (
            .O(N__19936),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1858 (
            .O(N__19933),
            .I(N__19930));
    InMux I__1857 (
            .O(N__19930),
            .I(N__19927));
    LocalMux I__1856 (
            .O(N__19927),
            .I(N__19924));
    Span4Mux_h I__1855 (
            .O(N__19924),
            .I(N__19921));
    Odrv4 I__1854 (
            .O(N__19921),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1853 (
            .O(N__19918),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1852 (
            .O(N__19915),
            .I(N__19912));
    InMux I__1851 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__1850 (
            .O(N__19909),
            .I(N__19906));
    Span4Mux_v I__1849 (
            .O(N__19906),
            .I(N__19903));
    Odrv4 I__1848 (
            .O(N__19903),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1847 (
            .O(N__19900),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__1846 (
            .O(N__19897),
            .I(N__19894));
    InMux I__1845 (
            .O(N__19894),
            .I(N__19891));
    LocalMux I__1844 (
            .O(N__19891),
            .I(N__19888));
    Span4Mux_h I__1843 (
            .O(N__19888),
            .I(N__19885));
    Odrv4 I__1842 (
            .O(N__19885),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1841 (
            .O(N__19882),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__1840 (
            .O(N__19879),
            .I(N__19876));
    InMux I__1839 (
            .O(N__19876),
            .I(N__19873));
    LocalMux I__1838 (
            .O(N__19873),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1837 (
            .O(N__19870),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__1836 (
            .O(N__19867),
            .I(N__19864));
    InMux I__1835 (
            .O(N__19864),
            .I(N__19861));
    LocalMux I__1834 (
            .O(N__19861),
            .I(N__19858));
    Span4Mux_h I__1833 (
            .O(N__19858),
            .I(N__19855));
    Odrv4 I__1832 (
            .O(N__19855),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1831 (
            .O(N__19852),
            .I(bfn_2_14_0_));
    CascadeMux I__1830 (
            .O(N__19849),
            .I(N__19846));
    InMux I__1829 (
            .O(N__19846),
            .I(N__19843));
    LocalMux I__1828 (
            .O(N__19843),
            .I(N__19840));
    Span4Mux_v I__1827 (
            .O(N__19840),
            .I(N__19837));
    Odrv4 I__1826 (
            .O(N__19837),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1825 (
            .O(N__19834),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1824 (
            .O(N__19831),
            .I(N__19828));
    InMux I__1823 (
            .O(N__19828),
            .I(N__19825));
    LocalMux I__1822 (
            .O(N__19825),
            .I(N__19822));
    Span4Mux_v I__1821 (
            .O(N__19822),
            .I(N__19819));
    Odrv4 I__1820 (
            .O(N__19819),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__1819 (
            .O(N__19816),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1818 (
            .O(N__19813),
            .I(N__19810));
    InMux I__1817 (
            .O(N__19810),
            .I(N__19807));
    LocalMux I__1816 (
            .O(N__19807),
            .I(N__19804));
    Span4Mux_h I__1815 (
            .O(N__19804),
            .I(N__19801));
    Span4Mux_s0_h I__1814 (
            .O(N__19801),
            .I(N__19798));
    Odrv4 I__1813 (
            .O(N__19798),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1812 (
            .O(N__19795),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1811 (
            .O(N__19792),
            .I(N__19789));
    InMux I__1810 (
            .O(N__19789),
            .I(N__19786));
    LocalMux I__1809 (
            .O(N__19786),
            .I(N__19783));
    Span4Mux_v I__1808 (
            .O(N__19783),
            .I(N__19780));
    Span4Mux_h I__1807 (
            .O(N__19780),
            .I(N__19777));
    Odrv4 I__1806 (
            .O(N__19777),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1805 (
            .O(N__19774),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__1804 (
            .O(N__19771),
            .I(N__19768));
    InMux I__1803 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__1802 (
            .O(N__19765),
            .I(N__19762));
    Span4Mux_v I__1801 (
            .O(N__19762),
            .I(N__19759));
    Span4Mux_h I__1800 (
            .O(N__19759),
            .I(N__19756));
    Odrv4 I__1799 (
            .O(N__19756),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1798 (
            .O(N__19753),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1797 (
            .O(N__19750),
            .I(N__19747));
    InMux I__1796 (
            .O(N__19747),
            .I(N__19744));
    LocalMux I__1795 (
            .O(N__19744),
            .I(N__19741));
    Span4Mux_h I__1794 (
            .O(N__19741),
            .I(N__19738));
    Odrv4 I__1793 (
            .O(N__19738),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1792 (
            .O(N__19735),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    InMux I__1791 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__1790 (
            .O(N__19729),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1789 (
            .O(N__19726),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    InMux I__1788 (
            .O(N__19723),
            .I(N__19720));
    LocalMux I__1787 (
            .O(N__19720),
            .I(N__19717));
    Odrv4 I__1786 (
            .O(N__19717),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1785 (
            .O(N__19714),
            .I(bfn_2_13_0_));
    CascadeMux I__1784 (
            .O(N__19711),
            .I(N__19708));
    InMux I__1783 (
            .O(N__19708),
            .I(N__19705));
    LocalMux I__1782 (
            .O(N__19705),
            .I(N__19702));
    Odrv4 I__1781 (
            .O(N__19702),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1780 (
            .O(N__19699),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1779 (
            .O(N__19696),
            .I(N__19693));
    InMux I__1778 (
            .O(N__19693),
            .I(N__19690));
    LocalMux I__1777 (
            .O(N__19690),
            .I(N__19687));
    Odrv4 I__1776 (
            .O(N__19687),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1775 (
            .O(N__19684),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__1774 (
            .O(N__19681),
            .I(N__19678));
    InMux I__1773 (
            .O(N__19678),
            .I(N__19675));
    LocalMux I__1772 (
            .O(N__19675),
            .I(N__19672));
    Span4Mux_h I__1771 (
            .O(N__19672),
            .I(N__19669));
    Odrv4 I__1770 (
            .O(N__19669),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1769 (
            .O(N__19666),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1768 (
            .O(N__19663),
            .I(N__19660));
    InMux I__1767 (
            .O(N__19660),
            .I(N__19657));
    LocalMux I__1766 (
            .O(N__19657),
            .I(N__19654));
    Span4Mux_h I__1765 (
            .O(N__19654),
            .I(N__19651));
    Odrv4 I__1764 (
            .O(N__19651),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__1763 (
            .O(N__19648),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1762 (
            .O(N__19645),
            .I(N__19642));
    InMux I__1761 (
            .O(N__19642),
            .I(N__19639));
    LocalMux I__1760 (
            .O(N__19639),
            .I(N__19636));
    Span4Mux_v I__1759 (
            .O(N__19636),
            .I(N__19633));
    Span4Mux_h I__1758 (
            .O(N__19633),
            .I(N__19630));
    Odrv4 I__1757 (
            .O(N__19630),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1756 (
            .O(N__19627),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1755 (
            .O(N__19624),
            .I(N__19621));
    InMux I__1754 (
            .O(N__19621),
            .I(N__19618));
    LocalMux I__1753 (
            .O(N__19618),
            .I(N__19615));
    Span4Mux_v I__1752 (
            .O(N__19615),
            .I(N__19612));
    Span4Mux_h I__1751 (
            .O(N__19612),
            .I(N__19609));
    Odrv4 I__1750 (
            .O(N__19609),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1749 (
            .O(N__19606),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1748 (
            .O(N__19603),
            .I(N__19600));
    InMux I__1747 (
            .O(N__19600),
            .I(N__19597));
    LocalMux I__1746 (
            .O(N__19597),
            .I(N__19594));
    Span4Mux_v I__1745 (
            .O(N__19594),
            .I(N__19591));
    Odrv4 I__1744 (
            .O(N__19591),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1743 (
            .O(N__19588),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1742 (
            .O(N__19585),
            .I(N__19582));
    InMux I__1741 (
            .O(N__19582),
            .I(N__19579));
    LocalMux I__1740 (
            .O(N__19579),
            .I(N__19576));
    Span4Mux_h I__1739 (
            .O(N__19576),
            .I(N__19573));
    Span4Mux_s0_h I__1738 (
            .O(N__19573),
            .I(N__19570));
    Odrv4 I__1737 (
            .O(N__19570),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1736 (
            .O(N__19567),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__1735 (
            .O(N__19564),
            .I(N__19561));
    InMux I__1734 (
            .O(N__19561),
            .I(N__19558));
    LocalMux I__1733 (
            .O(N__19558),
            .I(N__19555));
    Span4Mux_h I__1732 (
            .O(N__19555),
            .I(N__19552));
    Odrv4 I__1731 (
            .O(N__19552),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1730 (
            .O(N__19549),
            .I(bfn_2_12_0_));
    CascadeMux I__1729 (
            .O(N__19546),
            .I(N__19543));
    InMux I__1728 (
            .O(N__19543),
            .I(N__19540));
    LocalMux I__1727 (
            .O(N__19540),
            .I(N__19537));
    Span4Mux_h I__1726 (
            .O(N__19537),
            .I(N__19534));
    Odrv4 I__1725 (
            .O(N__19534),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1724 (
            .O(N__19531),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1723 (
            .O(N__19528),
            .I(N__19525));
    InMux I__1722 (
            .O(N__19525),
            .I(N__19522));
    LocalMux I__1721 (
            .O(N__19522),
            .I(N__19519));
    Span4Mux_h I__1720 (
            .O(N__19519),
            .I(N__19516));
    Span4Mux_s0_h I__1719 (
            .O(N__19516),
            .I(N__19513));
    Odrv4 I__1718 (
            .O(N__19513),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1717 (
            .O(N__19510),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__1716 (
            .O(N__19507),
            .I(N__19504));
    LocalMux I__1715 (
            .O(N__19504),
            .I(N__19501));
    Span4Mux_v I__1714 (
            .O(N__19501),
            .I(N__19498));
    Odrv4 I__1713 (
            .O(N__19498),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1712 (
            .O(N__19495),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1711 (
            .O(N__19492),
            .I(N__19489));
    LocalMux I__1710 (
            .O(N__19489),
            .I(N__19486));
    Span4Mux_v I__1709 (
            .O(N__19486),
            .I(N__19483));
    Odrv4 I__1708 (
            .O(N__19483),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1707 (
            .O(N__19480),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1706 (
            .O(N__19477),
            .I(N__19474));
    LocalMux I__1705 (
            .O(N__19474),
            .I(N__19471));
    Span4Mux_v I__1704 (
            .O(N__19471),
            .I(N__19468));
    Odrv4 I__1703 (
            .O(N__19468),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1702 (
            .O(N__19465),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1701 (
            .O(N__19462),
            .I(N__19459));
    LocalMux I__1700 (
            .O(N__19459),
            .I(N__19456));
    Span4Mux_v I__1699 (
            .O(N__19456),
            .I(N__19453));
    Odrv4 I__1698 (
            .O(N__19453),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__1697 (
            .O(N__19450),
            .I(N__19436));
    CascadeMux I__1696 (
            .O(N__19449),
            .I(N__19433));
    CascadeMux I__1695 (
            .O(N__19448),
            .I(N__19430));
    CascadeMux I__1694 (
            .O(N__19447),
            .I(N__19427));
    CascadeMux I__1693 (
            .O(N__19446),
            .I(N__19424));
    CascadeMux I__1692 (
            .O(N__19445),
            .I(N__19421));
    CascadeMux I__1691 (
            .O(N__19444),
            .I(N__19418));
    CascadeMux I__1690 (
            .O(N__19443),
            .I(N__19415));
    CascadeMux I__1689 (
            .O(N__19442),
            .I(N__19412));
    CascadeMux I__1688 (
            .O(N__19441),
            .I(N__19409));
    CascadeMux I__1687 (
            .O(N__19440),
            .I(N__19406));
    CascadeMux I__1686 (
            .O(N__19439),
            .I(N__19403));
    LocalMux I__1685 (
            .O(N__19436),
            .I(N__19400));
    InMux I__1684 (
            .O(N__19433),
            .I(N__19393));
    InMux I__1683 (
            .O(N__19430),
            .I(N__19393));
    InMux I__1682 (
            .O(N__19427),
            .I(N__19393));
    InMux I__1681 (
            .O(N__19424),
            .I(N__19384));
    InMux I__1680 (
            .O(N__19421),
            .I(N__19384));
    InMux I__1679 (
            .O(N__19418),
            .I(N__19384));
    InMux I__1678 (
            .O(N__19415),
            .I(N__19384));
    InMux I__1677 (
            .O(N__19412),
            .I(N__19379));
    InMux I__1676 (
            .O(N__19409),
            .I(N__19379));
    InMux I__1675 (
            .O(N__19406),
            .I(N__19374));
    InMux I__1674 (
            .O(N__19403),
            .I(N__19374));
    Odrv4 I__1673 (
            .O(N__19400),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1672 (
            .O(N__19393),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1671 (
            .O(N__19384),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1670 (
            .O(N__19379),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1669 (
            .O(N__19374),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1668 (
            .O(N__19363),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1667 (
            .O(N__19360),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1666 (
            .O(N__19357),
            .I(N__19354));
    LocalMux I__1665 (
            .O(N__19354),
            .I(un7_start_stop_0_a3));
    CascadeMux I__1664 (
            .O(N__19351),
            .I(N__19348));
    InMux I__1663 (
            .O(N__19348),
            .I(N__19345));
    LocalMux I__1662 (
            .O(N__19345),
            .I(N__19342));
    Span4Mux_h I__1661 (
            .O(N__19342),
            .I(N__19339));
    Odrv4 I__1660 (
            .O(N__19339),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1659 (
            .O(N__19336),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__1658 (
            .O(N__19333),
            .I(N__19330));
    LocalMux I__1657 (
            .O(N__19330),
            .I(N__19327));
    Span4Mux_v I__1656 (
            .O(N__19327),
            .I(N__19324));
    Odrv4 I__1655 (
            .O(N__19324),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1654 (
            .O(N__19321),
            .I(N__19318));
    InMux I__1653 (
            .O(N__19318),
            .I(N__19315));
    LocalMux I__1652 (
            .O(N__19315),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1651 (
            .O(N__19312),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__1650 (
            .O(N__19309),
            .I(N__19306));
    LocalMux I__1649 (
            .O(N__19306),
            .I(N__19303));
    Span4Mux_v I__1648 (
            .O(N__19303),
            .I(N__19300));
    Odrv4 I__1647 (
            .O(N__19300),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1646 (
            .O(N__19297),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__1645 (
            .O(N__19294),
            .I(N__19291));
    LocalMux I__1644 (
            .O(N__19291),
            .I(N__19288));
    Span4Mux_v I__1643 (
            .O(N__19288),
            .I(N__19285));
    Odrv4 I__1642 (
            .O(N__19285),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1641 (
            .O(N__19282),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1640 (
            .O(N__19279),
            .I(N__19276));
    LocalMux I__1639 (
            .O(N__19276),
            .I(N__19273));
    Span4Mux_v I__1638 (
            .O(N__19273),
            .I(N__19270));
    Odrv4 I__1637 (
            .O(N__19270),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1636 (
            .O(N__19267),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__1635 (
            .O(N__19264),
            .I(N__19261));
    LocalMux I__1634 (
            .O(N__19261),
            .I(N__19258));
    Span4Mux_v I__1633 (
            .O(N__19258),
            .I(N__19255));
    Odrv4 I__1632 (
            .O(N__19255),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1631 (
            .O(N__19252),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1630 (
            .O(N__19249),
            .I(N__19246));
    LocalMux I__1629 (
            .O(N__19246),
            .I(N__19243));
    Span4Mux_v I__1628 (
            .O(N__19243),
            .I(N__19240));
    Odrv4 I__1627 (
            .O(N__19240),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1626 (
            .O(N__19237),
            .I(bfn_1_12_0_));
    InMux I__1625 (
            .O(N__19234),
            .I(N__19231));
    LocalMux I__1624 (
            .O(N__19231),
            .I(N__19228));
    Span4Mux_v I__1623 (
            .O(N__19228),
            .I(N__19225));
    Odrv4 I__1622 (
            .O(N__19225),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1621 (
            .O(N__19222),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1620 (
            .O(N__19219),
            .I(N__19216));
    LocalMux I__1619 (
            .O(N__19216),
            .I(N__19213));
    Span4Mux_v I__1618 (
            .O(N__19213),
            .I(N__19210));
    Odrv4 I__1617 (
            .O(N__19210),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1616 (
            .O(N__19207),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1615 (
            .O(N__19204),
            .I(N__19201));
    LocalMux I__1614 (
            .O(N__19201),
            .I(N__19198));
    Span4Mux_v I__1613 (
            .O(N__19198),
            .I(N__19195));
    Odrv4 I__1612 (
            .O(N__19195),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1611 (
            .O(N__19192),
            .I(N__19189));
    LocalMux I__1610 (
            .O(N__19189),
            .I(N__19186));
    Span4Mux_v I__1609 (
            .O(N__19186),
            .I(N__19183));
    Odrv4 I__1608 (
            .O(N__19183),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1607 (
            .O(N__19180),
            .I(N__19177));
    InMux I__1606 (
            .O(N__19177),
            .I(N__19174));
    LocalMux I__1605 (
            .O(N__19174),
            .I(N__19171));
    Odrv4 I__1604 (
            .O(N__19171),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1603 (
            .O(N__19168),
            .I(N__19165));
    LocalMux I__1602 (
            .O(N__19165),
            .I(N__19162));
    Span4Mux_v I__1601 (
            .O(N__19162),
            .I(N__19159));
    Odrv4 I__1600 (
            .O(N__19159),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1599 (
            .O(N__19156),
            .I(N__19153));
    InMux I__1598 (
            .O(N__19153),
            .I(N__19150));
    LocalMux I__1597 (
            .O(N__19150),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1596 (
            .O(N__19147),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1595 (
            .O(N__19144),
            .I(N__19141));
    LocalMux I__1594 (
            .O(N__19141),
            .I(N__19138));
    Span4Mux_v I__1593 (
            .O(N__19138),
            .I(N__19135));
    Odrv4 I__1592 (
            .O(N__19135),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1591 (
            .O(N__19132),
            .I(N__19129));
    InMux I__1590 (
            .O(N__19129),
            .I(N__19126));
    LocalMux I__1589 (
            .O(N__19126),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1588 (
            .O(N__19123),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    IoInMux I__1587 (
            .O(N__19120),
            .I(N__19117));
    LocalMux I__1586 (
            .O(N__19117),
            .I(N__19114));
    Span4Mux_s3_v I__1585 (
            .O(N__19114),
            .I(N__19111));
    Span4Mux_h I__1584 (
            .O(N__19111),
            .I(N__19108));
    Sp12to4 I__1583 (
            .O(N__19108),
            .I(N__19105));
    Span12Mux_v I__1582 (
            .O(N__19105),
            .I(N__19102));
    Span12Mux_v I__1581 (
            .O(N__19102),
            .I(N__19099));
    Odrv12 I__1580 (
            .O(N__19099),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1579 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__1578 (
            .O(N__19093),
            .I(N__19090));
    IoSpan4Mux I__1577 (
            .O(N__19090),
            .I(N__19087));
    IoSpan4Mux I__1576 (
            .O(N__19087),
            .I(N__19084));
    Odrv4 I__1575 (
            .O(N__19084),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_16_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_27_0_));
    defparam IN_MUX_bfv_16_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_28_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_16_28_0_));
    defparam IN_MUX_bfv_16_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_29_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_16_29_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_27_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_13_27_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_17_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_27_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_17_27_0_));
    defparam IN_MUX_bfv_17_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_28_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_17_28_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_12_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_26_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_8_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_8_24_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_7_17_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19120),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19096),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__21124),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_161_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__46879),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__41269),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__40546),
            .CLKHFEN(N__40612),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__40478),
            .RGB2PWM(N__19957),
            .RGB1(rgb_g),
            .CURREN(N__40511),
            .RGB2(rgb_b),
            .RGB1PWM(N__19357),
            .RGB0PWM(N__49555),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__19204),
            .in2(_gnd_net_),
            .in3(N__19450),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__19192),
            .in2(N__19180),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__19168),
            .in2(N__19156),
            .in3(N__19147),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__19144),
            .in2(N__19132),
            .in3(N__19123),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__19333),
            .in2(N__19321),
            .in3(N__19312),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__19309),
            .in2(N__19439),
            .in3(N__19297),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__19294),
            .in2(N__19441),
            .in3(N__19282),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__19279),
            .in2(N__19440),
            .in3(N__19267),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19264),
            .in2(N__19442),
            .in3(N__19252),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__19249),
            .in2(N__19443),
            .in3(N__19237),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__19234),
            .in2(N__19447),
            .in3(N__19222),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__19219),
            .in2(N__19444),
            .in3(N__19207),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__19507),
            .in2(N__19448),
            .in3(N__19495),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__19492),
            .in2(N__19445),
            .in3(N__19480),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__19477),
            .in2(N__19449),
            .in3(N__19465),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__19462),
            .in2(N__19446),
            .in3(N__19363),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19360),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_24_0  (
            .in0(N__43339),
            .in1(N__40317),
            .in2(_gnd_net_),
            .in3(N__42376),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_0_a3_LC_1_29_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_0_a3_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_0_a3_LC_1_29_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un7_start_stop_0_a3_LC_1_29_0  (
            .in0(N__49554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44812),
            .lcout(un7_start_stop_0_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__39916),
            .in2(N__20235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__37064),
            .in2(N__19351),
            .in3(N__19336),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__37006),
            .in2(N__19681),
            .in3(N__19666),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__36946),
            .in2(N__19663),
            .in3(N__19648),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__36910),
            .in2(N__19645),
            .in3(N__19627),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__36820),
            .in2(N__19624),
            .in3(N__19606),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__37582),
            .in2(N__19603),
            .in3(N__19588),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__37534),
            .in2(N__19585),
            .in3(N__19567),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__37471),
            .in2(N__19564),
            .in3(N__19549),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__37414),
            .in2(N__19546),
            .in3(N__19531),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__37341),
            .in2(N__19528),
            .in3(N__19510),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__37267),
            .in2(N__19813),
            .in3(N__19795),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__37207),
            .in2(N__19792),
            .in3(N__19774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__37153),
            .in2(N__19771),
            .in3(N__19753),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__38029),
            .in2(N__19750),
            .in3(N__19735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__19732),
            .in2(N__37983),
            .in3(N__19726),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__19723),
            .in2(N__37926),
            .in3(N__19714),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__37876),
            .in2(N__19711),
            .in3(N__19699),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__37822),
            .in2(N__19696),
            .in3(N__19684),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__37762),
            .in2(N__19948),
            .in3(N__19936),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__37699),
            .in2(N__19933),
            .in3(N__19918),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__37645),
            .in2(N__19915),
            .in3(N__19900),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__38503),
            .in2(N__19897),
            .in3(N__19882),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__38437),
            .in2(N__19879),
            .in3(N__19870),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__38384),
            .in2(N__19867),
            .in3(N__19852),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__38329),
            .in2(N__19849),
            .in3(N__19834),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__38257),
            .in2(N__19831),
            .in3(N__19816),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__38213),
            .in2(N__20068),
            .in3(N__20053),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__38156),
            .in2(N__20050),
            .in3(N__20038),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__38092),
            .in2(N__20035),
            .in3(N__20020),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_14_6  (
            .in0(N__20017),
            .in1(N__38708),
            .in2(N__20008),
            .in3(N__19993),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_0 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_0  (
            .in0(N__20672),
            .in1(N__38730),
            .in2(N__19990),
            .in3(N__20377),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(),
            .sr(N__49513));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_15_1 .LUT_INIT=16'b1100010011000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_2_15_1  (
            .in0(N__38729),
            .in1(N__19981),
            .in2(N__20426),
            .in3(N__20675),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(),
            .sr(N__49513));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_15_5 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_2_15_5  (
            .in0(N__38728),
            .in1(N__20674),
            .in2(N__20425),
            .in3(N__19972),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(),
            .sr(N__49513));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_6 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_6  (
            .in0(N__20673),
            .in1(N__38731),
            .in2(N__19966),
            .in3(N__20378),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(),
            .sr(N__49513));
    defparam \phase_controller_inst1.N_39_i_i_LC_2_30_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_39_i_i_LC_2_30_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_39_i_i_LC_2_30_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.N_39_i_i_LC_2_30_7  (
            .in0(_gnd_net_),
            .in1(N__44811),
            .in2(_gnd_net_),
            .in3(N__49553),
            .lcout(N_39_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_11_0 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_3_11_0  (
            .in0(N__20422),
            .in1(N__38803),
            .in2(N__20687),
            .in3(N__20134),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50013),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_11_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_3_11_1  (
            .in0(N__20128),
            .in1(N__20655),
            .in2(_gnd_net_),
            .in3(N__20423),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50013),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_11_7 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_3_11_7  (
            .in0(N__38802),
            .in1(N__20656),
            .in2(N__20122),
            .in3(N__20424),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50013),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_12_0 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_3_12_0  (
            .in0(N__20420),
            .in1(N__38779),
            .in2(N__20690),
            .in3(N__20113),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50005),
            .ce(),
            .sr(N__49495));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2  (
            .in0(N__20419),
            .in1(_gnd_net_),
            .in2(N__20689),
            .in3(N__20104),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50005),
            .ce(),
            .sr(N__49495));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_12_3 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_3_12_3  (
            .in0(N__38777),
            .in1(N__20660),
            .in2(N__20098),
            .in3(N__20421),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50005),
            .ce(),
            .sr(N__49495));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_12_4 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_12_4  (
            .in0(N__20418),
            .in1(N__38778),
            .in2(N__20688),
            .in3(N__20089),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50005),
            .ce(),
            .sr(N__49495));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_13_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_3_13_2  (
            .in0(N__38782),
            .in1(N__20403),
            .in2(N__20083),
            .in3(N__20652),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_13_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_3_13_3  (
            .in0(N__20650),
            .in1(N__38784),
            .in2(N__20434),
            .in3(N__20074),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_13_4 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_3_13_4  (
            .in0(N__38783),
            .in1(N__20404),
            .in2(N__20203),
            .in3(N__20653),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_13_5 .LUT_INIT=16'b1100111111001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_3_13_5  (
            .in0(N__20649),
            .in1(N__20194),
            .in2(N__20436),
            .in3(N__38786),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_13_7 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_3_13_7  (
            .in0(N__20651),
            .in1(N__38785),
            .in2(N__20435),
            .in3(N__20188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_14_0 .LUT_INIT=16'b1101110111001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_3_14_0  (
            .in0(N__20398),
            .in1(N__20182),
            .in2(N__20691),
            .in3(N__38736),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_1 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_1  (
            .in0(N__38733),
            .in1(N__20400),
            .in2(N__20176),
            .in3(N__20685),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_14_2 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_3_14_2  (
            .in0(N__20399),
            .in1(N__38735),
            .in2(N__20692),
            .in3(N__20167),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_14_5 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_3_14_5  (
            .in0(N__38734),
            .in1(N__20401),
            .in2(N__20161),
            .in3(N__20686),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_7 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_7  (
            .in0(N__38732),
            .in1(N__20678),
            .in2(N__20152),
            .in3(N__20402),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_3_15_2 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_3_15_2  (
            .in0(N__20677),
            .in1(N__38738),
            .in2(N__20428),
            .in3(N__20140),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49509));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_15_4 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_3_15_4  (
            .in0(N__20676),
            .in1(N__38737),
            .in2(N__20427),
            .in3(N__20266),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49509));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_0  (
            .in0(N__38212),
            .in1(N__38383),
            .in2(N__38264),
            .in3(N__38333),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_2  (
            .in0(N__20260),
            .in1(N__20242),
            .in2(N__20254),
            .in3(N__20734),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_4  (
            .in0(N__37703),
            .in1(N__38699),
            .in2(N__38447),
            .in3(N__37763),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_16_6  (
            .in0(N__38040),
            .in1(N__37223),
            .in2(N__37427),
            .in3(N__37976),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_7  (
            .in0(N__38100),
            .in1(N__37287),
            .in2(N__20245),
            .in3(N__20275),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_3_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_3_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_3_17_2  (
            .in0(N__37925),
            .in1(N__37830),
            .in2(N__37656),
            .in3(N__37878),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_3_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_3_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_3_17_6  (
            .in0(N__37283),
            .in1(N__37340),
            .in2(N__37170),
            .in3(N__37975),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_11_5 .LUT_INIT=16'b0011110000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_4_11_5  (
            .in0(N__20623),
            .in1(N__39915),
            .in2(N__20236),
            .in3(N__20433),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50006),
            .ce(),
            .sr(N__49487));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_4_12_0 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_4_12_0  (
            .in0(N__20429),
            .in1(N__38792),
            .in2(N__20670),
            .in3(N__20212),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(),
            .sr(N__49492));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_1 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_1  (
            .in0(N__38790),
            .in1(N__20615),
            .in2(N__20515),
            .in3(N__20431),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(),
            .sr(N__49492));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_12_4 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_4_12_4  (
            .in0(N__20430),
            .in1(N__38793),
            .in2(N__20671),
            .in3(N__20503),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(),
            .sr(N__49492));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_12_7 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_4_12_7  (
            .in0(N__38791),
            .in1(N__20616),
            .in2(N__20494),
            .in3(N__20432),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(),
            .sr(N__49492));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_4_13_1 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_4_13_1  (
            .in0(N__20654),
            .in1(N__38781),
            .in2(N__20479),
            .in3(N__20417),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49987),
            .ce(),
            .sr(N__49496));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_14_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_4_14_3  (
            .in0(N__20597),
            .in1(N__38799),
            .in2(N__20437),
            .in3(N__20464),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49974),
            .ce(),
            .sr(N__49500));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_4_15_5 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_4_15_5  (
            .in0(N__38800),
            .in1(N__20598),
            .in2(N__20452),
            .in3(N__20385),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49963),
            .ce(),
            .sr(N__49504));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__37163),
            .in2(_gnd_net_),
            .in3(N__37330),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_16_2  (
            .in0(N__37536),
            .in1(N__37592),
            .in2(N__36848),
            .in3(N__37475),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_16_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_16_3  (
            .in0(N__36965),
            .in1(N__37025),
            .in2(N__20269),
            .in3(N__36915),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_16_4  (
            .in0(N__38152),
            .in1(N__38504),
            .in2(N__20737),
            .in3(N__20728),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_16_6  (
            .in0(N__37924),
            .in1(N__37823),
            .in2(N__37655),
            .in3(N__37877),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_0  (
            .in0(N__38036),
            .in1(N__37224),
            .in2(N__37434),
            .in3(N__38157),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_17_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__38337),
            .in2(_gnd_net_),
            .in3(N__37704),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_17_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_17_2  (
            .in0(N__38448),
            .in1(N__37764),
            .in2(N__20722),
            .in3(N__20521),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_3  (
            .in0(N__38511),
            .in1(N__38780),
            .in2(N__20719),
            .in3(N__20716),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_4  (
            .in0(N__20710),
            .in1(N__20701),
            .in2(N__20695),
            .in3(N__20767),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_17_7  (
            .in0(N__38220),
            .in1(N__38093),
            .in2(N__38271),
            .in3(N__38388),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_5_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_5_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_5_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_5_8_1  (
            .in0(N__26726),
            .in1(N__26707),
            .in2(_gnd_net_),
            .in3(N__30226),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50019),
            .ce(N__29275),
            .sr(N__49463));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_5_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_5_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_5_8_7  (
            .in0(N__27007),
            .in1(N__26963),
            .in2(_gnd_net_),
            .in3(N__30227),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50019),
            .ce(N__29275),
            .sr(N__49463));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_5_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_5_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_5_9_0  (
            .in0(N__30219),
            .in1(N__25994),
            .in2(_gnd_net_),
            .in3(N__26601),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_5_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_5_9_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_5_9_2  (
            .in0(N__20794),
            .in1(N__25819),
            .in2(N__23164),
            .in3(N__27001),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_5_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_5_9_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_5_9_3  (
            .in0(N__26727),
            .in1(_gnd_net_),
            .in2(N__20755),
            .in3(N__26705),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_5_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_5_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_5_9_5  (
            .in0(N__20817),
            .in1(N__21565),
            .in2(_gnd_net_),
            .in3(N__30221),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_5_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_5_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_5_9_6  (
            .in0(N__30220),
            .in1(N__27002),
            .in2(_gnd_net_),
            .in3(N__26967),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_5_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_5_10_3 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_5_10_3  (
            .in0(N__20778),
            .in1(N__23085),
            .in2(N__23119),
            .in3(N__20751),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_5_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_5_10_6 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_5_10_6  (
            .in0(N__23118),
            .in1(N__20752),
            .in2(N__23086),
            .in3(N__20779),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_5_10_7  (
            .in0(N__30225),
            .in1(N__20813),
            .in2(_gnd_net_),
            .in3(N__21563),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50007),
            .ce(N__29274),
            .sr(N__49477));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_5_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_5_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_5_11_4  (
            .in0(N__27081),
            .in1(N__27053),
            .in2(_gnd_net_),
            .in3(N__30246),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49998),
            .ce(N__29256),
            .sr(N__49483));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_5_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_5_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_5_11_5  (
            .in0(N__30245),
            .in1(N__24900),
            .in2(_gnd_net_),
            .in3(N__24876),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49998),
            .ce(N__29256),
            .sr(N__49483));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_5_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_5_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_5_12_0  (
            .in0(N__27231),
            .in1(N__30247),
            .in2(_gnd_net_),
            .in3(N__27208),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49988),
            .ce(N__29267),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_13_3  (
            .in0(N__26162),
            .in1(N__26141),
            .in2(_gnd_net_),
            .in3(N__30241),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_5_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_5_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_5_13_5  (
            .in0(N__24899),
            .in1(N__24875),
            .in2(_gnd_net_),
            .in3(N__30242),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_5_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_5_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_5_14_1  (
            .in0(N__27230),
            .in1(N__27206),
            .in2(_gnd_net_),
            .in3(N__30244),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_5_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_5_15_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_5_15_3  (
            .in0(N__27080),
            .in1(N__27057),
            .in2(_gnd_net_),
            .in3(N__30243),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_5_17_0 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_5_17_0  (
            .in0(N__37035),
            .in1(N__37080),
            .in2(N__39942),
            .in3(N__36975),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_5_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_5_17_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_5_17_1  (
            .in0(N__20761),
            .in1(N__37482),
            .in2(N__20770),
            .in3(N__36849),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_5_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_5_17_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_5_17_6  (
            .in0(N__36914),
            .in1(N__37535),
            .in2(_gnd_net_),
            .in3(N__37593),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_7_7_0  (
            .in0(N__26914),
            .in1(N__26930),
            .in2(_gnd_net_),
            .in3(N__30319),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50014),
            .ce(N__29235),
            .sr(N__49438));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_7_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_7_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_7_8_1  (
            .in0(N__26068),
            .in1(N__26593),
            .in2(N__21564),
            .in3(N__26912),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_7_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_7_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_7_8_6  (
            .in0(N__30368),
            .in1(N__20821),
            .in2(_gnd_net_),
            .in3(N__21559),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50008),
            .ce(N__30102),
            .sr(N__49446));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_9_0  (
            .in0(N__26615),
            .in1(N__26519),
            .in2(N__28636),
            .in3(N__29494),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_7_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_7_9_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_7_9_1  (
            .in0(N__24827),
            .in1(_gnd_net_),
            .in2(N__20797),
            .in3(N__30613),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21423),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49999),
            .ce(N__22645),
            .sr(N__49455));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21399),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49999),
            .ce(N__22645),
            .sr(N__49455));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_9_6  (
            .in0(N__26616),
            .in1(N__26645),
            .in2(_gnd_net_),
            .in3(N__30302),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_10_0  (
            .in0(N__22573),
            .in1(N__21419),
            .in2(_gnd_net_),
            .in3(N__20785),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_10_1  (
            .in0(N__22569),
            .in1(N__21395),
            .in2(_gnd_net_),
            .in3(N__20782),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_10_2  (
            .in0(N__22574),
            .in1(N__21376),
            .in2(_gnd_net_),
            .in3(N__20848),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_10_3  (
            .in0(N__22570),
            .in1(N__21354),
            .in2(_gnd_net_),
            .in3(N__20845),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_10_4  (
            .in0(N__22575),
            .in1(N__21332),
            .in2(_gnd_net_),
            .in3(N__20842),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_10_5  (
            .in0(N__22571),
            .in1(N__21306),
            .in2(_gnd_net_),
            .in3(N__20839),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_10_6  (
            .in0(N__22576),
            .in1(N__21286),
            .in2(_gnd_net_),
            .in3(N__20836),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_10_7  (
            .in0(N__22572),
            .in1(N__21268),
            .in2(_gnd_net_),
            .in3(N__20833),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__49989),
            .ce(N__22410),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_11_0  (
            .in0(N__22564),
            .in1(N__21641),
            .in2(_gnd_net_),
            .in3(N__20830),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_11_1  (
            .in0(N__22568),
            .in1(N__21608),
            .in2(_gnd_net_),
            .in3(N__20827),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_11_2  (
            .in0(N__22561),
            .in1(N__21582),
            .in2(_gnd_net_),
            .in3(N__20824),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_11_3  (
            .in0(N__22565),
            .in1(N__21526),
            .in2(_gnd_net_),
            .in3(N__20875),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_11_4  (
            .in0(N__22562),
            .in1(N__21504),
            .in2(_gnd_net_),
            .in3(N__20872),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_11_5  (
            .in0(N__22566),
            .in1(N__21482),
            .in2(_gnd_net_),
            .in3(N__20869),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_11_6  (
            .in0(N__22563),
            .in1(N__21460),
            .in2(_gnd_net_),
            .in3(N__20866),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_11_7  (
            .in0(N__22567),
            .in1(N__21442),
            .in2(_gnd_net_),
            .in3(N__20863),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49975),
            .ce(N__22411),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_12_0  (
            .in0(N__22529),
            .in1(N__21857),
            .in2(_gnd_net_),
            .in3(N__20860),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_12_1  (
            .in0(N__22548),
            .in1(N__21827),
            .in2(_gnd_net_),
            .in3(N__20857),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_12_2  (
            .in0(N__22530),
            .in1(N__21801),
            .in2(_gnd_net_),
            .in3(N__20854),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_12_3  (
            .in0(N__22549),
            .in1(N__21781),
            .in2(_gnd_net_),
            .in3(N__20851),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_12_4  (
            .in0(N__22531),
            .in1(N__21759),
            .in2(_gnd_net_),
            .in3(N__20902),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_12_5  (
            .in0(N__22550),
            .in1(N__21737),
            .in2(_gnd_net_),
            .in3(N__20899),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_12_6  (
            .in0(N__22532),
            .in1(N__21715),
            .in2(_gnd_net_),
            .in3(N__20896),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_12_7  (
            .in0(N__22551),
            .in1(N__21697),
            .in2(_gnd_net_),
            .in3(N__20893),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49964),
            .ce(N__22409),
            .sr(N__49478));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_13_0  (
            .in0(N__22542),
            .in1(N__21671),
            .in2(_gnd_net_),
            .in3(N__20890),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_13_1  (
            .in0(N__22546),
            .in1(N__21995),
            .in2(_gnd_net_),
            .in3(N__20887),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_13_2  (
            .in0(N__22543),
            .in1(N__21957),
            .in2(_gnd_net_),
            .in3(N__20884),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_13_3  (
            .in0(N__22547),
            .in1(N__21923),
            .in2(_gnd_net_),
            .in3(N__20881),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_13_4  (
            .in0(N__22544),
            .in1(N__21973),
            .in2(_gnd_net_),
            .in3(N__20878),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_13_5  (
            .in0(N__21937),
            .in1(N__22545),
            .in2(_gnd_net_),
            .in3(N__20932),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49955),
            .ce(N__22399),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__20929),
            .in2(_gnd_net_),
            .in3(N__21898),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__21892),
            .in2(_gnd_net_),
            .in3(N__20923),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__21883),
            .in2(_gnd_net_),
            .in3(N__20920),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__21874),
            .in2(_gnd_net_),
            .in3(N__20917),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__22078),
            .in2(_gnd_net_),
            .in3(N__20914),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__22069),
            .in2(_gnd_net_),
            .in3(N__20911),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__22060),
            .in2(_gnd_net_),
            .in3(N__20908),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__22051),
            .in2(_gnd_net_),
            .in3(N__20905),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49489));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__22042),
            .in2(_gnd_net_),
            .in3(N__20959),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__22033),
            .in2(_gnd_net_),
            .in3(N__20956),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__22024),
            .in2(_gnd_net_),
            .in3(N__20953),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__22015),
            .in2(_gnd_net_),
            .in3(N__20950),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__22006),
            .in2(_gnd_net_),
            .in3(N__20947),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_7_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__22150),
            .in2(_gnd_net_),
            .in3(N__20944),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_7_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__22141),
            .in2(_gnd_net_),
            .in3(N__20941),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_7_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_7_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__22132),
            .in2(_gnd_net_),
            .in3(N__20938),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__49939),
            .ce(),
            .sr(N__49493));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_7_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__22123),
            .in2(_gnd_net_),
            .in3(N__20935),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_7_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__22114),
            .in2(_gnd_net_),
            .in3(N__20986),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_7_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_7_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__22105),
            .in2(_gnd_net_),
            .in3(N__20983),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_7_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__22096),
            .in2(_gnd_net_),
            .in3(N__20980),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_7_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_7_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__22087),
            .in2(_gnd_net_),
            .in3(N__20977),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_7_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_7_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__22225),
            .in2(_gnd_net_),
            .in3(N__20974),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_7_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_7_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_7_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__22216),
            .in2(_gnd_net_),
            .in3(N__20971),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_7_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_7_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_7_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__22207),
            .in2(_gnd_net_),
            .in3(N__20968),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49497));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_7_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_7_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__22198),
            .in2(_gnd_net_),
            .in3(N__20965),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_7_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_7_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__22189),
            .in2(_gnd_net_),
            .in3(N__20962),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_7_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_7_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_7_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__22180),
            .in2(_gnd_net_),
            .in3(N__21097),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_7_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_7_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_7_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__22171),
            .in2(_gnd_net_),
            .in3(N__21094),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_7_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_7_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_7_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__22162),
            .in2(_gnd_net_),
            .in3(N__21091),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_7_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_7_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_7_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__22300),
            .in2(_gnd_net_),
            .in3(N__21088),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_7_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_7_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_7_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__22255),
            .in2(_gnd_net_),
            .in3(N__21085),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_7_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_7_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__22267),
            .in2(_gnd_net_),
            .in3(N__21082),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49501));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21066),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49505));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_7_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_7_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21048),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49505));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_7_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_7_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_7_19_5  (
            .in0(N__21030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(),
            .sr(N__49510));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21006),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21186),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_7_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_7_24_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_7_24_2  (
            .in0(N__22756),
            .in1(N__21144),
            .in2(_gnd_net_),
            .in3(N__21164),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_7_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_7_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_7_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21143),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_7_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_7_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_7_25_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_7_25_0  (
            .in0(N__24054),
            .in1(N__42463),
            .in2(N__22762),
            .in3(N__21165),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.timer_s1.running_LC_7_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_7_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_7_25_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_7_25_7  (
            .in0(N__21166),
            .in1(N__22760),
            .in2(_gnd_net_),
            .in3(N__21145),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_26_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_7_26_7  (
            .in0(_gnd_net_),
            .in1(N__21163),
            .in2(_gnd_net_),
            .in3(N__21142),
            .lcout(\current_shift_inst.timer_s1.N_161_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_8_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_8_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_8_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22355),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(),
            .sr(N__49415));
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22356),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(),
            .sr(N__49415));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_6_4  (
            .in0(N__26072),
            .in1(N__26030),
            .in2(_gnd_net_),
            .in3(N__30330),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_8_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_8_6_6 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_8_6_6  (
            .in0(N__23061),
            .in1(N__21250),
            .in2(N__23035),
            .in3(N__21235),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_6_7  (
            .in0(N__30329),
            .in1(N__26934),
            .in2(_gnd_net_),
            .in3(N__26911),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_7_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_7_1  (
            .in0(N__21249),
            .in1(N__23028),
            .in2(N__23062),
            .in3(N__21234),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_8_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_8_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_8_7_2  (
            .in0(N__26860),
            .in1(N__26820),
            .in2(_gnd_net_),
            .in3(N__30303),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_8_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_8_7_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_8_7_3  (
            .in0(N__30304),
            .in1(_gnd_net_),
            .in2(N__21238),
            .in3(N__26861),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50009),
            .ce(N__29215),
            .sr(N__49430));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_8_7_6  (
            .in0(N__26001),
            .in1(N__26594),
            .in2(_gnd_net_),
            .in3(N__30305),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50009),
            .ce(N__29215),
            .sr(N__49430));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_8_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_8_8_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_8_8_0  (
            .in0(N__21220),
            .in1(N__22983),
            .in2(N__21211),
            .in3(N__23001),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_8_1  (
            .in0(N__26792),
            .in1(N__26754),
            .in2(_gnd_net_),
            .in3(N__30356),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_8_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_8_8_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_8_8_2  (
            .in0(N__30357),
            .in1(_gnd_net_),
            .in2(N__21223),
            .in3(N__26793),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50000),
            .ce(N__29255),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_8_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_8_8_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_8_8_4  (
            .in0(N__21219),
            .in1(N__22982),
            .in2(N__21210),
            .in3(N__23000),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__21374),
            .in2(N__21424),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__21353),
            .in2(N__21403),
            .in3(N__21379),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__21375),
            .in2(N__21333),
            .in3(N__21361),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__21305),
            .in2(N__21358),
            .in3(N__21337),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__21284),
            .in2(N__21334),
            .in3(N__21313),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__21266),
            .in2(N__21310),
            .in3(N__21289),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__21285),
            .in2(N__21649),
            .in3(N__21271),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__21267),
            .in2(N__21619),
            .in3(N__21253),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49990),
            .ce(N__22644),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__21581),
            .in2(N__21648),
            .in3(N__21622),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__21524),
            .in2(N__21615),
            .in3(N__21589),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__21503),
            .in2(N__21586),
            .in3(N__21529),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__21525),
            .in2(N__21483),
            .in3(N__21511),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__21458),
            .in2(N__21508),
            .in3(N__21487),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__21440),
            .in2(N__21484),
            .in3(N__21463),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__21459),
            .in2(N__21865),
            .in3(N__21445),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__21441),
            .in2(N__21835),
            .in3(N__21427),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49976),
            .ce(N__22643),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__21800),
            .in2(N__21864),
            .in3(N__21838),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__21779),
            .in2(N__21834),
            .in3(N__21808),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__21758),
            .in2(N__21805),
            .in3(N__21784),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__21780),
            .in2(N__21738),
            .in3(N__21766),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__21713),
            .in2(N__21763),
            .in3(N__21742),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__21695),
            .in2(N__21739),
            .in3(N__21718),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__21714),
            .in2(N__21679),
            .in3(N__21700),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__21696),
            .in2(N__22000),
            .in3(N__21682),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49965),
            .ce(N__22642),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__21956),
            .in2(N__21678),
            .in3(N__21652),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49956),
            .ce(N__22629),
            .sr(N__49470));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__21996),
            .in2(N__21924),
            .in3(N__21976),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49956),
            .ce(N__22629),
            .sr(N__49470));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__21972),
            .in2(N__21961),
            .in3(N__21940),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49956),
            .ce(N__22629),
            .sr(N__49470));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__21936),
            .in2(N__21925),
            .in3(N__21904),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49956),
            .ce(N__22629),
            .sr(N__49470));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21901),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__22629),
            .sr(N__49470));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__23302),
            .in2(N__23290),
            .in3(N__23288),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__23380),
            .in2(_gnd_net_),
            .in3(N__21886),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__23251),
            .in2(_gnd_net_),
            .in3(N__21877),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_13_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__23257),
            .in2(_gnd_net_),
            .in3(N__21868),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_13_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__23368),
            .in2(_gnd_net_),
            .in3(N__22072),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_13_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__23362),
            .in2(_gnd_net_),
            .in3(N__22063),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__23356),
            .in2(_gnd_net_),
            .in3(N__22054),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__22423),
            .in2(_gnd_net_),
            .in3(N__22045),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__23320),
            .in2(_gnd_net_),
            .in3(N__22036),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__23269),
            .in2(_gnd_net_),
            .in3(N__22027),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__23350),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__23263),
            .in2(_gnd_net_),
            .in3(N__22009),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_14_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__23338),
            .in2(_gnd_net_),
            .in3(N__22153),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__23344),
            .in2(_gnd_net_),
            .in3(N__22144),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_8_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_8_14_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__23326),
            .in2(_gnd_net_),
            .in3(N__22135),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_8_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_8_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__23404),
            .in2(_gnd_net_),
            .in3(N__22126),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_8_15_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__23374),
            .in2(_gnd_net_),
            .in3(N__22117),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_8_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__22441),
            .in2(_gnd_net_),
            .in3(N__22108),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_8_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__22288),
            .in2(_gnd_net_),
            .in3(N__22099),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_8_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__22432),
            .in2(_gnd_net_),
            .in3(N__22090),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_8_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__23332),
            .in2(_gnd_net_),
            .in3(N__22081),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_8_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__22276),
            .in2(_gnd_net_),
            .in3(N__22219),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_8_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__22249),
            .in2(_gnd_net_),
            .in3(N__22210),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_8_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__22240),
            .in2(_gnd_net_),
            .in3(N__22201),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_8_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__22231),
            .in2(_gnd_net_),
            .in3(N__22192),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_8_16_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__22582),
            .in2(_gnd_net_),
            .in3(N__22183),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_8_16_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23398),
            .in3(N__22174),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_8_16_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__22282),
            .in2(_gnd_net_),
            .in3(N__22165),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_8_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__25243),
            .in2(_gnd_net_),
            .in3(N__22156),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_8_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_8_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__23314),
            .in2(_gnd_net_),
            .in3(N__22294),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_8_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(_gnd_net_),
            .in3(N__22291),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_16_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_16_7  (
            .in0(N__25376),
            .in1(N__25009),
            .in2(_gnd_net_),
            .in3(N__27988),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_8_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_8_17_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_8_17_0  (
            .in0(N__25352),
            .in1(N__28090),
            .in2(_gnd_net_),
            .in3(N__25390),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_1  (
            .in0(N__27928),
            .in1(N__25156),
            .in2(_gnd_net_),
            .in3(N__25347),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_8_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_8_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4  (
            .in0(N__25348),
            .in1(N__27913),
            .in2(_gnd_net_),
            .in3(N__25144),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_17_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_17_5  (
            .in0(N__25132),
            .in1(N__27883),
            .in2(_gnd_net_),
            .in3(N__25349),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_17_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_17_6  (
            .in0(N__25350),
            .in1(N__28138),
            .in2(_gnd_net_),
            .in3(N__25120),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_17_7 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_17_7  (
            .in0(N__25108),
            .in1(N__25351),
            .in2(_gnd_net_),
            .in3(N__28123),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_18_0  (
            .in0(N__22333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_18_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_18_1  (
            .in0(N__28003),
            .in1(N__25024),
            .in2(_gnd_net_),
            .in3(N__25294),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_18_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_18_4  (
            .in0(N__25295),
            .in1(N__25180),
            .in2(_gnd_net_),
            .in3(N__27958),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_8_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_8_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_8_18_5  (
            .in0(N__35551),
            .in1(N__25758),
            .in2(N__35237),
            .in3(N__28459),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_18_7  (
            .in0(N__32778),
            .in1(N__31952),
            .in2(_gnd_net_),
            .in3(N__31989),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_19_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_19_0  (
            .in0(N__27595),
            .in1(N__24949),
            .in2(_gnd_net_),
            .in3(N__25293),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_19_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_19_1  (
            .in0(N__22317),
            .in1(N__22334),
            .in2(_gnd_net_),
            .in3(N__22362),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_199_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_19_2 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_8_19_2  (
            .in0(N__22363),
            .in1(_gnd_net_),
            .in2(N__22339),
            .in3(N__22318),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49506));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_19_4  (
            .in0(N__22335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22316),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_198_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_19_6 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_8_19_6  (
            .in0(N__28975),
            .in1(N__48554),
            .in2(_gnd_net_),
            .in3(N__48516),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32248),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_20_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__35602),
            .in2(N__22597),
            .in3(N__32953),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32183),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__32881),
            .sr(N__49511));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_20_4  (
            .in0(N__32211),
            .in1(N__40616),
            .in2(_gnd_net_),
            .in3(N__22594),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_20_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_20_5  (
            .in0(N__40617),
            .in1(_gnd_net_),
            .in2(N__22588),
            .in3(N__27501),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_8_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_8_20_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_8_20_6  (
            .in0(N__32489),
            .in1(N__32777),
            .in2(_gnd_net_),
            .in3(N__32469),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_8_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_8_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32488),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_8_21_0  (
            .in0(N__22921),
            .in1(N__32970),
            .in2(_gnd_net_),
            .in3(N__22585),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_8_21_1  (
            .in0(N__22917),
            .in1(N__32898),
            .in2(_gnd_net_),
            .in3(N__22672),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_8_21_2  (
            .in0(N__22922),
            .in1(N__23618),
            .in2(_gnd_net_),
            .in3(N__22669),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_8_21_3  (
            .in0(N__22918),
            .in1(N__23588),
            .in2(_gnd_net_),
            .in3(N__22666),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_8_21_4  (
            .in0(N__22923),
            .in1(N__23568),
            .in2(_gnd_net_),
            .in3(N__22663),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_8_21_5  (
            .in0(N__22919),
            .in1(N__23544),
            .in2(_gnd_net_),
            .in3(N__22660),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_8_21_6  (
            .in0(N__22924),
            .in1(N__23521),
            .in2(_gnd_net_),
            .in3(N__22657),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_8_21_7  (
            .in0(N__22920),
            .in1(N__23503),
            .in2(_gnd_net_),
            .in3(N__22654),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49894),
            .ce(N__22798),
            .sr(N__49515));
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_8_22_0  (
            .in0(N__22912),
            .in1(N__23477),
            .in2(_gnd_net_),
            .in3(N__22651),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_8_22_1  (
            .in0(N__22916),
            .in1(N__23447),
            .in2(_gnd_net_),
            .in3(N__22648),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_8_22_2  (
            .in0(N__22909),
            .in1(N__23832),
            .in2(_gnd_net_),
            .in3(N__22699),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_8_22_3  (
            .in0(N__22913),
            .in1(N__23809),
            .in2(_gnd_net_),
            .in3(N__22696),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_8_22_4  (
            .in0(N__22910),
            .in1(N__23790),
            .in2(_gnd_net_),
            .in3(N__22693),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_8_22_5  (
            .in0(N__22914),
            .in1(N__23765),
            .in2(_gnd_net_),
            .in3(N__22690),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_8_22_6  (
            .in0(N__22911),
            .in1(N__23743),
            .in2(_gnd_net_),
            .in3(N__22687),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_8_22_7  (
            .in0(N__22915),
            .in1(N__23725),
            .in2(_gnd_net_),
            .in3(N__22684),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49887),
            .ce(N__22797),
            .sr(N__49519));
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_8_23_0  (
            .in0(N__22881),
            .in1(N__23702),
            .in2(_gnd_net_),
            .in3(N__22681),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_8_23_1  (
            .in0(N__22885),
            .in1(N__23669),
            .in2(_gnd_net_),
            .in3(N__22678),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_8_23_2  (
            .in0(N__22882),
            .in1(N__23643),
            .in2(_gnd_net_),
            .in3(N__22675),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_8_23_3  (
            .in0(N__22886),
            .in1(N__24031),
            .in2(_gnd_net_),
            .in3(N__22726),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_8_23_4  (
            .in0(N__22883),
            .in1(N__24012),
            .in2(_gnd_net_),
            .in3(N__22723),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_8_23_5  (
            .in0(N__22887),
            .in1(N__23987),
            .in2(_gnd_net_),
            .in3(N__22720),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_8_23_6  (
            .in0(N__22884),
            .in1(N__23965),
            .in2(_gnd_net_),
            .in3(N__22717),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_8_23_7  (
            .in0(N__22888),
            .in1(N__23947),
            .in2(_gnd_net_),
            .in3(N__22714),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49882),
            .ce(N__22784),
            .sr(N__49522));
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_8_24_0  (
            .in0(N__22877),
            .in1(N__23924),
            .in2(_gnd_net_),
            .in3(N__22711),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_8_24_1  (
            .in0(N__22889),
            .in1(N__23894),
            .in2(_gnd_net_),
            .in3(N__22708),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_8_24_2  (
            .in0(N__22878),
            .in1(N__23856),
            .in2(_gnd_net_),
            .in3(N__22705),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_8_24_3  (
            .in0(N__22890),
            .in1(N__24090),
            .in2(_gnd_net_),
            .in3(N__22702),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_8_24_4  (
            .in0(N__22879),
            .in1(N__23869),
            .in2(_gnd_net_),
            .in3(N__22927),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_8_24_5  (
            .in0(N__24103),
            .in1(N__22880),
            .in2(_gnd_net_),
            .in3(N__22801),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(N__22783),
            .sr(N__49524));
    defparam \current_shift_inst.start_timer_s1_LC_8_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_8_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_8_25_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_8_25_4  (
            .in0(N__24047),
            .in1(N__22761),
            .in2(_gnd_net_),
            .in3(N__42461),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(),
            .sr(N__49526));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_9_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_9_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_9_6_3  (
            .in0(N__26452),
            .in1(N__26409),
            .in2(_gnd_net_),
            .in3(N__30328),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_9_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_9_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__24193),
            .in2(N__25849),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_7_1  (
            .in0(N__29186),
            .in1(N__24172),
            .in2(_gnd_net_),
            .in3(N__22738),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_7_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_7_2  (
            .in0(N__29190),
            .in1(N__24151),
            .in2(N__24205),
            .in3(N__22735),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_7_3  (
            .in0(N__29187),
            .in1(N__24124),
            .in2(_gnd_net_),
            .in3(N__22732),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_7_4  (
            .in0(N__29191),
            .in1(N__24370),
            .in2(_gnd_net_),
            .in3(N__22729),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_7_5  (
            .in0(N__29188),
            .in1(N__24349),
            .in2(_gnd_net_),
            .in3(N__22954),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_7_6  (
            .in0(N__29192),
            .in1(N__24331),
            .in2(_gnd_net_),
            .in3(N__22951),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_7_7  (
            .in0(N__29189),
            .in1(N__24310),
            .in2(_gnd_net_),
            .in3(N__22948),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50001),
            .ce(),
            .sr(N__49423));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_8_0  (
            .in0(N__29124),
            .in1(N__24292),
            .in2(_gnd_net_),
            .in3(N__22945),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_8_1  (
            .in0(N__29117),
            .in1(N__24274),
            .in2(_gnd_net_),
            .in3(N__22942),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_8_2  (
            .in0(N__29121),
            .in1(N__24256),
            .in2(_gnd_net_),
            .in3(N__22939),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_8_3  (
            .in0(N__29118),
            .in1(N__24232),
            .in2(_gnd_net_),
            .in3(N__22936),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_8_4  (
            .in0(N__29122),
            .in1(N__24538),
            .in2(_gnd_net_),
            .in3(N__22933),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_8_5  (
            .in0(N__29119),
            .in1(N__24502),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_8_6  (
            .in0(N__29123),
            .in1(N__24472),
            .in2(_gnd_net_),
            .in3(N__23065),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_8_7  (
            .in0(N__29120),
            .in1(N__23060),
            .in2(_gnd_net_),
            .in3(N__23038),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49991),
            .ce(),
            .sr(N__49431));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_9_0  (
            .in0(N__29193),
            .in1(N__23027),
            .in2(_gnd_net_),
            .in3(N__23005),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_9_1  (
            .in0(N__29239),
            .in1(N__23002),
            .in2(_gnd_net_),
            .in3(N__22987),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_9_2  (
            .in0(N__29194),
            .in1(N__22984),
            .in2(_gnd_net_),
            .in3(N__22969),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_9_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_9_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_9_9_3  (
            .in0(N__29240),
            .in1(N__25931),
            .in2(_gnd_net_),
            .in3(N__22966),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_9_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_9_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_9_9_4  (
            .in0(N__29195),
            .in1(N__25952),
            .in2(_gnd_net_),
            .in3(N__22963),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_9_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_9_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_9_9_5  (
            .in0(N__29241),
            .in1(N__24692),
            .in2(_gnd_net_),
            .in3(N__22960),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_9_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_9_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_9_9_6  (
            .in0(N__29196),
            .in1(N__24710),
            .in2(_gnd_net_),
            .in3(N__22957),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_9_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_9_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_9_9_7  (
            .in0(N__29242),
            .in1(N__23195),
            .in2(_gnd_net_),
            .in3(N__23137),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49977),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_9_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_9_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_9_10_0  (
            .in0(N__29223),
            .in1(N__23233),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_9_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_9_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_9_10_1  (
            .in0(N__29236),
            .in1(N__24574),
            .in2(_gnd_net_),
            .in3(N__23131),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_9_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_9_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_9_10_2  (
            .in0(N__29224),
            .in1(N__24591),
            .in2(_gnd_net_),
            .in3(N__23128),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_9_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_9_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_9_10_3  (
            .in0(N__29237),
            .in1(N__26210),
            .in2(_gnd_net_),
            .in3(N__23125),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_9_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_9_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_9_10_4  (
            .in0(N__29225),
            .in1(N__26231),
            .in2(_gnd_net_),
            .in3(N__23122),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_9_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_9_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_9_10_5  (
            .in0(N__29238),
            .in1(N__23108),
            .in2(_gnd_net_),
            .in3(N__23092),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_9_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_9_10_6  (
            .in0(N__29226),
            .in1(N__23081),
            .in2(_gnd_net_),
            .in3(N__23089),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49966),
            .ce(),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_9_11_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_9_11_0  (
            .in0(N__23242),
            .in1(N__23232),
            .in2(N__23218),
            .in3(N__23197),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_11_1  (
            .in0(N__26321),
            .in1(N__26298),
            .in2(_gnd_net_),
            .in3(N__30526),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(elapsed_time_ns_1_RNI25DN9_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_11_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_9_11_2  (
            .in0(N__30527),
            .in1(_gnd_net_),
            .in2(N__23245),
            .in3(N__26322),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49957),
            .ce(N__29266),
            .sr(N__49457));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_11_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_11_4  (
            .in0(N__23241),
            .in1(N__23231),
            .in2(N__23217),
            .in3(N__23196),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_1  (
            .in0(N__26791),
            .in1(N__26686),
            .in2(N__26865),
            .in3(N__29447),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_12_2  (
            .in0(N__23149),
            .in1(N__23143),
            .in2(N__23179),
            .in3(N__23176),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_9_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_9_12_3 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__28995),
            .in2(N__48571),
            .in3(N__48517),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_201_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_12_4  (
            .in0(N__30659),
            .in1(N__24856),
            .in2(N__26131),
            .in3(N__27040),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_12_6  (
            .in0(N__26380),
            .in1(N__26342),
            .in2(_gnd_net_),
            .in3(N__30346),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_12_7  (
            .in0(N__27187),
            .in1(N__27267),
            .in2(N__26480),
            .in3(N__26320),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_9_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_9_13_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_9_13_0  (
            .in0(N__24934),
            .in1(N__27868),
            .in2(_gnd_net_),
            .in3(N__25358),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_13_1  (
            .in0(N__25360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_9_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_9_13_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_9_13_2  (
            .in0(N__24790),
            .in1(N__27721),
            .in2(_gnd_net_),
            .in3(N__25356),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_9_13_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23293),
            .in3(N__23289),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49471));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25357),
            .lcout(\current_shift_inst.N_1306_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_9_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_9_13_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_9_13_7  (
            .in0(N__25359),
            .in1(N__27850),
            .in2(_gnd_net_),
            .in3(N__24922),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_9_14_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_9_14_0  (
            .in0(N__25367),
            .in1(N__25081),
            .in2(_gnd_net_),
            .in3(N__27811),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_9_14_1 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_9_14_1  (
            .in0(N__24988),
            .in1(N__25363),
            .in2(_gnd_net_),
            .in3(N__27667),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_9_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_9_14_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_9_14_2  (
            .in0(N__25362),
            .in1(N__27682),
            .in2(_gnd_net_),
            .in3(N__24997),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_9_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_9_14_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_9_14_3  (
            .in0(N__27703),
            .in1(N__24781),
            .in2(_gnd_net_),
            .in3(N__25361),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_9_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_9_14_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_9_14_4  (
            .in0(N__25368),
            .in1(N__28030),
            .in2(_gnd_net_),
            .in3(N__25036),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_9_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_9_14_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_9_14_5  (
            .in0(N__27652),
            .in1(N__24976),
            .in2(_gnd_net_),
            .in3(N__25364),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_9_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_9_14_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_9_14_6  (
            .in0(N__25365),
            .in1(N__24967),
            .in2(_gnd_net_),
            .in3(N__27634),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_9_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_9_14_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_9_14_7  (
            .in0(N__27616),
            .in1(N__24958),
            .in2(_gnd_net_),
            .in3(N__25366),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_9_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_9_15_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_9_15_0  (
            .in0(N__24910),
            .in1(N__27826),
            .in2(_gnd_net_),
            .in3(N__25369),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_9_15_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_9_15_1  (
            .in0(N__25371),
            .in1(N__25063),
            .in2(_gnd_net_),
            .in3(N__27778),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_9_15_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_9_15_2  (
            .in0(N__27796),
            .in1(N__25072),
            .in2(_gnd_net_),
            .in3(N__25370),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_3  (
            .in0(N__25374),
            .in1(N__27943),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_9_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_9_15_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_9_15_4  (
            .in0(N__27760),
            .in1(N__25054),
            .in2(_gnd_net_),
            .in3(N__25372),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_9_15_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_9_15_5  (
            .in0(N__25373),
            .in1(N__27739),
            .in2(_gnd_net_),
            .in3(N__25045),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_9_15_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_9_15_6  (
            .in0(N__28108),
            .in1(N__25093),
            .in2(_gnd_net_),
            .in3(N__25375),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__32584),
            .in2(N__32215),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__40732),
            .in2(N__32617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__25549),
            .in2(N__40755),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__40736),
            .in2(N__25486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__25561),
            .in2(N__40756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__40740),
            .in2(N__27448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__23389),
            .in2(N__40757),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__40744),
            .in2(N__27427),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__40728),
            .in2(N__31834),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__32263),
            .in2(N__40754),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__40716),
            .in2(N__25198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__23416),
            .in2(N__40751),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__40720),
            .in2(N__25471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__25222),
            .in2(N__40752),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__40724),
            .in2(N__25216),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__25588),
            .in2(N__40753),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__40659),
            .in2(N__25462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__25231),
            .in2(N__40712),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__40663),
            .in2(N__25663),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__25414),
            .in2(N__40713),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__40667),
            .in2(N__25645),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__25789),
            .in2(N__40714),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__40671),
            .in2(N__25408),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__25189),
            .in2(N__40715),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__40618),
            .in2(N__25576),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25537),
            .in2(N__40656),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__40622),
            .in2(N__25681),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25435),
            .in2(N__40657),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__40626),
            .in2(N__25453),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__25516),
            .in2(N__40658),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__40630),
            .in2(N__25444),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__35595),
            .in2(_gnd_net_),
            .in3(N__23422),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_9_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_9_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__32969),
            .in2(N__23619),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__32897),
            .in2(N__23595),
            .in3(N__23419),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_9_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(N__23620),
            .in3(N__23599),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__23540),
            .in2(N__23596),
            .in3(N__23572),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_9_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__23519),
            .in2(N__23569),
            .in3(N__23548),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__23501),
            .in2(N__23545),
            .in3(N__23524),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_9_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__23520),
            .in2(N__23485),
            .in3(N__23506),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_9_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__23502),
            .in2(N__23452),
            .in3(N__23488),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49895),
            .ce(N__32880),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__23828),
            .in2(N__23481),
            .in3(N__23455),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__23807),
            .in2(N__23451),
            .in3(N__23425),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__23786),
            .in2(N__23833),
            .in3(N__23812),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__23808),
            .in2(N__23766),
            .in3(N__23794),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__23741),
            .in2(N__23791),
            .in3(N__23770),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__23723),
            .in2(N__23767),
            .in3(N__23746),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__23742),
            .in2(N__23707),
            .in3(N__23728),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_9_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__23724),
            .in2(N__23676),
            .in3(N__23710),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49888),
            .ce(N__32879),
            .sr(N__49512));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_9_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__23639),
            .in2(N__23706),
            .in3(N__23680),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_9_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__24029),
            .in2(N__23677),
            .in3(N__23647),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_9_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__24008),
            .in2(N__23644),
            .in3(N__23623),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_9_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__24030),
            .in2(N__23988),
            .in3(N__24016),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_9_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__23963),
            .in2(N__24013),
            .in3(N__23992),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_9_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_9_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__23945),
            .in2(N__23989),
            .in3(N__23968),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_9_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_9_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_9_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__23964),
            .in2(N__23929),
            .in3(N__23950),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_9_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_9_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_9_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__23946),
            .in2(N__23899),
            .in3(N__23932),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49883),
            .ce(N__32877),
            .sr(N__49516));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_9_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_9_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__23852),
            .in2(N__23928),
            .in3(N__23902),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49879),
            .ce(N__32876),
            .sr(N__49520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_9_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__24086),
            .in2(N__23898),
            .in3(N__23872),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49879),
            .ce(N__32876),
            .sr(N__49520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_9_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_9_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__23868),
            .in2(N__23857),
            .in3(N__23836),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49879),
            .ce(N__32876),
            .sr(N__49520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_9_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_9_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__24102),
            .in2(N__24091),
            .in3(N__24070),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49879),
            .ce(N__32876),
            .sr(N__49520));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_9_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_9_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24067),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31348),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_9_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_9_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_9_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42462),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(),
            .sr(N__49525));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_10_5_7  (
            .in0(N__28668),
            .in1(N__28650),
            .in2(_gnd_net_),
            .in3(N__30432),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50002),
            .ce(N__29219),
            .sr(N__49397));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_10_6_0  (
            .in0(N__30421),
            .in1(N__26555),
            .in2(_gnd_net_),
            .in3(N__26538),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49992),
            .ce(N__29246),
            .sr(N__49403));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_1  (
            .in0(N__26460),
            .in1(N__26405),
            .in2(_gnd_net_),
            .in3(N__30423),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49992),
            .ce(N__29246),
            .sr(N__49403));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_10_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_10_6_3  (
            .in0(N__26034),
            .in1(N__26076),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49992),
            .ce(N__29246),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28994),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_10_7_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_10_7_1  (
            .in0(N__37125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28577),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_7_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_7_2  (
            .in0(N__28575),
            .in1(N__25872),
            .in2(_gnd_net_),
            .in3(N__37124),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_10_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24208),
            .in3(N__25860),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_10_7_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_10_7_4  (
            .in0(N__28576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28547),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_7_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24196),
            .in3(N__28603),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_10_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_10_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__24187),
            .in2(N__25882),
            .in3(N__25838),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_10_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_10_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__24181),
            .in2(N__24160),
            .in3(N__24171),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_10_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_10_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__24139),
            .in2(N__24655),
            .in3(N__24150),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_10_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_10_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__24133),
            .in2(N__24112),
            .in3(N__24123),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_10_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_10_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__24379),
            .in2(N__24358),
            .in3(N__24369),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_10_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_10_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__24337),
            .in2(N__24604),
            .in3(N__24348),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_10_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_10_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__26185),
            .in2(N__24319),
            .in3(N__24330),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_10_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_10_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__24298),
            .in2(N__29290),
            .in3(N__24309),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_10_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_10_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_10_9_0  (
            .in0(N__24291),
            .in1(N__24280),
            .in2(N__25978),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_10_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_10_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__24262),
            .in2(N__25798),
            .in3(N__24273),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_10_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__25969),
            .in2(N__24244),
            .in3(N__24255),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_10_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_10_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__29299),
            .in2(N__24220),
            .in3(N__24231),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_10_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_10_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__24553),
            .in2(N__24526),
            .in3(N__24537),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_10_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_10_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__24514),
            .in2(N__24490),
            .in3(N__24501),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_10_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_10_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__24481),
            .in2(N__24460),
            .in3(N__24471),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_10_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_10_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__24451),
            .in2(N__24439),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_10_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__24424),
            .in2(N__24412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_10_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_10_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__25915),
            .in2(N__25963),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_10_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_10_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__24676),
            .in2(N__24745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_10_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_10_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__24397),
            .in2(N__24388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_10_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_10_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__24559),
            .in2(N__24616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_10_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_10_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__26194),
            .in2(N__26245),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_10_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_10_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__24643),
            .in2(N__24631),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24619),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0  (
            .in0(N__24573),
            .in1(N__24754),
            .in2(N__24769),
            .in3(N__24590),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_11_1  (
            .in0(N__30501),
            .in1(N__26285),
            .in2(_gnd_net_),
            .in3(N__26256),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(elapsed_time_ns_1_RNII43T9_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_10_11_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_10_11_2  (
            .in0(N__26286),
            .in1(_gnd_net_),
            .in2(N__24607),
            .in3(N__30504),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49942),
            .ce(N__29265),
            .sr(N__49441));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_11_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_11_3  (
            .in0(N__24753),
            .in1(N__24768),
            .in2(N__24592),
            .in3(N__24572),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_10_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_10_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_10_11_4  (
            .in0(N__24836),
            .in1(N__24801),
            .in2(_gnd_net_),
            .in3(N__30500),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(elapsed_time_ns_1_RNI58DN9_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_11_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_10_11_5  (
            .in0(N__30503),
            .in1(_gnd_net_),
            .in2(N__24772),
            .in3(N__24837),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49942),
            .ce(N__29265),
            .sr(N__49441));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_10_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_10_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_10_11_6  (
            .in0(N__30668),
            .in1(N__30639),
            .in2(_gnd_net_),
            .in3(N__30499),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(elapsed_time_ns_1_RNI47DN9_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_10_11_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_10_11_7  (
            .in0(N__30502),
            .in1(_gnd_net_),
            .in2(N__24757),
            .in3(N__30669),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49942),
            .ce(N__29265),
            .sr(N__49441));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_12_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_12_0  (
            .in0(N__24694),
            .in1(N__24664),
            .in2(N__24730),
            .in3(N__24714),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_10_12_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_10_12_1  (
            .in0(N__24663),
            .in1(N__24729),
            .in2(N__24715),
            .in3(N__24693),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_12_4  (
            .in0(N__27281),
            .in1(N__27252),
            .in2(_gnd_net_),
            .in3(N__30429),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_10_12_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_10_12_5  (
            .in0(N__30430),
            .in1(_gnd_net_),
            .in2(N__24667),
            .in3(N__27282),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49931),
            .ce(N__29254),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_10_12_6  (
            .in0(N__26652),
            .in1(N__26628),
            .in2(_gnd_net_),
            .in3(N__30431),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49931),
            .ce(N__29254),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_10_13_0  (
            .in0(N__30426),
            .in1(N__26169),
            .in2(_gnd_net_),
            .in3(N__26143),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__30097),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_13_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_10_13_1  (
            .in0(N__27116),
            .in1(_gnd_net_),
            .in2(N__27157),
            .in3(N__30427),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__30097),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_10_13_5  (
            .in0(N__24901),
            .in1(N__24877),
            .in2(_gnd_net_),
            .in3(N__30428),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__30097),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_10_13_6  (
            .in0(N__30425),
            .in1(N__24838),
            .in2(_gnd_net_),
            .in3(N__24805),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__30097),
            .sr(N__49458));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_10_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_10_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__25498),
            .in2(N__27535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_10_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__32822),
            .in2(N__32926),
            .in3(N__32596),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_10_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_10_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_10_14_2  (
            .in0(N__32597),
            .in1(N__34719),
            .in2(N__30931),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_10_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__31000),
            .in2(N__34869),
            .in3(N__24784),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_10_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__34723),
            .in2(N__25531),
            .in3(N__24775),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_10_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__25399),
            .in2(N__34870),
            .in3(N__24991),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_10_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__34727),
            .in2(N__25429),
            .in3(N__24979),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_10_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_10_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__31744),
            .in2(N__34871),
            .in3(N__24970),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_10_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__34731),
            .in2(N__27487),
            .in3(N__24961),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_10_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__32347),
            .in2(N__34872),
            .in3(N__24952),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_10_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__34735),
            .in2(N__27547),
            .in3(N__24937),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_10_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__25600),
            .in2(N__34873),
            .in3(N__24925),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_10_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__34739),
            .in2(N__27436),
            .in3(N__24913),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_10_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__25609),
            .in2(N__34874),
            .in3(N__24904),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_10_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__34743),
            .in2(N__27358),
            .in3(N__25075),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_10_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__26947),
            .in2(N__34875),
            .in3(N__25066),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_10_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__34977),
            .in2(N__27295),
            .in3(N__25057),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_10_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__27577),
            .in2(N__35136),
            .in3(N__25048),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_10_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__34981),
            .in2(N__25696),
            .in3(N__25039),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_10_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__27583),
            .in2(N__35137),
            .in3(N__25027),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_10_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_10_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__34985),
            .in2(N__27304),
            .in3(N__25012),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_10_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_10_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__27346),
            .in2(N__35138),
            .in3(N__25000),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_10_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_10_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__34989),
            .in2(N__27367),
            .in3(N__25168),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_10_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_10_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__27571),
            .in2(N__35139),
            .in3(N__25159),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_10_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_10_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__35000),
            .in2(N__27565),
            .in3(N__25147),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_10_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_10_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__25777),
            .in2(N__35143),
            .in3(N__25135),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_10_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_10_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__35004),
            .in2(N__25729),
            .in3(N__25123),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_10_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_10_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__27556),
            .in2(N__35144),
            .in3(N__25111),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_10_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_10_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__35008),
            .in2(N__25714),
            .in3(N__25096),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_10_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__25768),
            .in2(N__35145),
            .in3(N__25084),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_10_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_10_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__35012),
            .in2(N__25207),
            .in3(N__25381),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_10_17_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_10_17_7  (
            .in0(N__32320),
            .in1(N__28069),
            .in2(N__25378),
            .in3(N__25246),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_18_0  (
            .in0(N__32783),
            .in1(N__31358),
            .in2(_gnd_net_),
            .in3(N__31401),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_18_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_18_1  (
            .in0(N__25630),
            .in1(N__35534),
            .in2(N__28387),
            .in3(N__35184),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_18_2  (
            .in0(N__32781),
            .in1(N__25629),
            .in2(_gnd_net_),
            .in3(N__28383),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_3  (
            .in0(N__31079),
            .in1(N__32782),
            .in2(_gnd_net_),
            .in3(N__30908),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_4  (
            .in0(N__35185),
            .in1(N__35535),
            .in2(N__32598),
            .in3(N__32542),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_18_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_18_5  (
            .in0(N__32138),
            .in1(N__32779),
            .in2(_gnd_net_),
            .in3(N__32113),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_18_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_18_6  (
            .in0(N__32784),
            .in1(N__34637),
            .in2(_gnd_net_),
            .in3(N__35283),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_18_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_18_7  (
            .in0(N__31684),
            .in1(N__32780),
            .in2(_gnd_net_),
            .in3(N__31715),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_19_0  (
            .in0(N__32761),
            .in1(N__30854),
            .in2(_gnd_net_),
            .in3(N__30809),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_19_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_19_1  (
            .in0(N__31302),
            .in1(N__35574),
            .in2(_gnd_net_),
            .in3(N__31269),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_10_19_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_10_19_2  (
            .in0(N__35576),
            .in1(N__35148),
            .in2(N__28254),
            .in3(N__27474),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_10_19_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__32541),
            .in2(_gnd_net_),
            .in3(N__35575),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_19_4  (
            .in0(N__35573),
            .in1(N__28856),
            .in2(_gnd_net_),
            .in3(N__28818),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_19_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_19_5  (
            .in0(N__35149),
            .in1(N__35577),
            .in2(N__31956),
            .in3(N__31985),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_19_6  (
            .in0(N__32762),
            .in1(N__31628),
            .in2(_gnd_net_),
            .in3(N__31599),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_19_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_19_7  (
            .in0(N__27411),
            .in1(N__32763),
            .in2(_gnd_net_),
            .in3(N__28518),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_10_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_10_20_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_10_20_0  (
            .in0(N__27473),
            .in1(N__35580),
            .in2(N__28255),
            .in3(N__35076),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_20_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_20_1  (
            .in0(N__31850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_20_2  (
            .in0(N__35552),
            .in1(N__31523),
            .in2(_gnd_net_),
            .in3(N__31557),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_20_3  (
            .in0(N__35579),
            .in1(N__31222),
            .in2(N__35192),
            .in3(N__31200),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32286),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_20_5  (
            .in0(N__35578),
            .in1(N__28770),
            .in2(_gnd_net_),
            .in3(N__28741),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31760),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_10_20_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_10_20_7  (
            .in0(N__25507),
            .in1(N__35553),
            .in2(_gnd_net_),
            .in3(N__32952),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_21_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_21_0  (
            .in0(N__28299),
            .in1(N__35583),
            .in2(N__35193),
            .in3(N__27329),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_21_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_21_1  (
            .in0(N__32743),
            .in1(N__30972),
            .in2(_gnd_net_),
            .in3(N__30948),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27469),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30971),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31942),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31457),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_21_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_21_6  (
            .in0(N__31227),
            .in1(N__32744),
            .in2(N__31199),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_21_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__31226),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_22_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_22_0  (
            .in0(N__32708),
            .in1(N__31475),
            .in2(_gnd_net_),
            .in3(N__31430),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32129),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31705),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25622),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_22_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_22_4  (
            .in0(N__25623),
            .in1(N__35582),
            .in2(N__28382),
            .in3(N__35197),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_10_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_10_22_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_10_22_5  (
            .in0(N__35581),
            .in1(N__32490),
            .in2(N__35238),
            .in3(N__32462),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_22_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_22_6  (
            .in0(N__32709),
            .in1(N__31142),
            .in2(_gnd_net_),
            .in3(N__31103),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31141),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32369),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_23_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_23_1  (
            .in0(N__32788),
            .in1(N__32023),
            .in2(_gnd_net_),
            .in3(N__32052),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27385),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30751),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31619),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27322),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_10_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_10_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35266),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_10_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_10_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30844),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_24_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_24_0  (
            .in0(N__35198),
            .in1(N__35604),
            .in2(N__30768),
            .in3(N__30729),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_24_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_24_1  (
            .in0(N__35603),
            .in1(N__25745),
            .in2(_gnd_net_),
            .in3(N__28445),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_24_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_24_2  (
            .in0(N__32785),
            .in1(N__30761),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_10_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_10_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31286),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28837),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25744),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_24_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_24_6  (
            .in0(N__32786),
            .in1(N__27330),
            .in2(_gnd_net_),
            .in3(N__28284),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_10_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_10_24_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_10_24_7  (
            .in0(N__32787),
            .in1(N__32376),
            .in2(_gnd_net_),
            .in3(N__32411),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32030),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_10_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_10_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28768),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_25_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_25_2  (
            .in0(N__35242),
            .in1(N__35606),
            .in2(N__31527),
            .in3(N__31550),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_25_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_25_3  (
            .in0(N__35609),
            .in1(N__35241),
            .in2(N__28740),
            .in3(N__28769),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_25_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_25_4  (
            .in0(N__35243),
            .in1(N__35607),
            .in2(N__28455),
            .in3(N__25759),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_10_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_10_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31519),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_25_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_25_6  (
            .in0(N__35239),
            .in1(N__35608),
            .in2(N__31268),
            .in3(N__31301),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_25_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_25_7  (
            .in0(N__35605),
            .in1(N__35240),
            .in2(N__27407),
            .in3(N__28511),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_11_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_11_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_11_6_0  (
            .in0(N__28669),
            .in1(N__28646),
            .in2(_gnd_net_),
            .in3(N__30420),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_11_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_11_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_11_6_4  (
            .in0(N__26559),
            .in1(N__26537),
            .in2(_gnd_net_),
            .in3(N__30419),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_7_2 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_11_7_2  (
            .in0(N__25873),
            .in1(N__28605),
            .in2(N__28584),
            .in3(N__28554),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49968),
            .ce(),
            .sr(N__49404));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37126),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49968),
            .ce(),
            .sr(N__49404));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_7_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_7_7  (
            .in0(N__28604),
            .in1(N__25861),
            .in2(N__25848),
            .in3(N__29149),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49968),
            .ce(),
            .sr(N__49404));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_11_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_11_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_11_8_0  (
            .in0(N__27151),
            .in1(N__28945),
            .in2(N__26389),
            .in3(N__28898),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_11_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_11_8_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_11_8_1  (
            .in0(N__26284),
            .in1(N__26459),
            .in2(N__25822),
            .in3(N__25807),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__29384),
            .in2(_gnd_net_),
            .in3(N__29351),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_11_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_11_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_11_8_4  (
            .in0(N__30493),
            .in1(N__28920),
            .in2(_gnd_net_),
            .in3(N__28946),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_5  (
            .in0(N__28947),
            .in1(_gnd_net_),
            .in2(N__25801),
            .in3(N__30497),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__29247),
            .sr(N__49409));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_6  (
            .in0(N__26387),
            .in1(_gnd_net_),
            .in2(N__30548),
            .in3(N__26349),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__29247),
            .sr(N__49409));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_7  (
            .in0(N__30557),
            .in1(N__27121),
            .in2(_gnd_net_),
            .in3(N__27152),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__29247),
            .sr(N__49409));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_11_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_11_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_11_9_0  (
            .in0(N__25954),
            .in1(N__25932),
            .in2(N__25906),
            .in3(N__25891),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_9_1  (
            .in0(N__25890),
            .in1(N__25953),
            .in2(N__25936),
            .in3(N__25902),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_11_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_11_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_11_9_2  (
            .in0(N__26489),
            .in1(N__26502),
            .in2(_gnd_net_),
            .in3(N__30437),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_11_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_11_9_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_11_9_3  (
            .in0(N__30440),
            .in1(_gnd_net_),
            .in2(N__25909),
            .in3(N__26490),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__29252),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_11_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_11_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_11_9_4  (
            .in0(N__29462),
            .in1(N__29430),
            .in2(_gnd_net_),
            .in3(N__30438),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_11_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_11_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_11_9_5  (
            .in0(N__30439),
            .in1(_gnd_net_),
            .in2(N__25894),
            .in3(N__29463),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__29252),
            .sr(N__49416));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_11_9_6  (
            .in0(N__29507),
            .in1(N__29539),
            .in2(_gnd_net_),
            .in3(N__30441),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__29252),
            .sr(N__49416));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_0  (
            .in0(N__26233),
            .in1(N__26211),
            .in2(N__26101),
            .in3(N__26086),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_10_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_10_1  (
            .in0(N__26085),
            .in1(N__26232),
            .in2(N__26215),
            .in3(N__26097),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_10_3  (
            .in0(N__30550),
            .in1(N__29360),
            .in2(_gnd_net_),
            .in3(N__29331),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_10_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_11_10_4  (
            .in0(N__29361),
            .in1(_gnd_net_),
            .in2(N__26188),
            .in3(N__30553),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__29248),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_11_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_11_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_11_10_5  (
            .in0(N__30552),
            .in1(N__26173),
            .in2(_gnd_net_),
            .in3(N__26142),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__29248),
            .sr(N__49424));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_11_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_11_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_11_10_6  (
            .in0(N__30617),
            .in1(N__30573),
            .in2(_gnd_net_),
            .in3(N__30549),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_11_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_11_10_7  (
            .in0(N__30551),
            .in1(_gnd_net_),
            .in2(N__26089),
            .in3(N__30618),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__29248),
            .sr(N__49424));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_11_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_11_11_0  (
            .in0(N__26077),
            .in1(_gnd_net_),
            .in2(N__30558),
            .in3(N__26038),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_11_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_11_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_11_11_1  (
            .in0(N__26008),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__30534),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_11_11_2  (
            .in0(N__30529),
            .in1(N__26563),
            .in2(_gnd_net_),
            .in3(N__26539),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_11_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_11_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_11_11_3  (
            .in0(N__26506),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(N__30535),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_11_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_11_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_11_11_4  (
            .in0(N__30530),
            .in1(N__26461),
            .in2(_gnd_net_),
            .in3(N__26416),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_11_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_11_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_11_11_5  (
            .in0(N__26388),
            .in1(N__26350),
            .in2(_gnd_net_),
            .in3(N__30537),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_11_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_11_11_6  (
            .in0(N__30528),
            .in1(N__26326),
            .in2(_gnd_net_),
            .in3(N__26302),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_11_11_7  (
            .in0(N__26287),
            .in1(N__26257),
            .in2(_gnd_net_),
            .in3(N__30536),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(N__30103),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_12_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_12_0  (
            .in0(N__33663),
            .in1(N__33636),
            .in2(N__26809),
            .in3(N__26875),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_12_1  (
            .in0(N__26874),
            .in1(N__33664),
            .in2(N__33640),
            .in3(N__26805),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_11_12_2  (
            .in0(N__26941),
            .in1(N__26913),
            .in2(_gnd_net_),
            .in3(N__30324),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(N__30101),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_11_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_11_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_11_12_3  (
            .in0(N__30323),
            .in1(N__26866),
            .in2(_gnd_net_),
            .in3(N__26830),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(N__30101),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_13_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_13_0  (
            .in0(N__33586),
            .in1(N__33609),
            .in2(N__26668),
            .in3(N__26743),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_11_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_11_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_11_13_1  (
            .in0(N__26742),
            .in1(N__33585),
            .in2(N__33613),
            .in3(N__26664),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_11_13_2  (
            .in0(N__30325),
            .in1(N__26797),
            .in2(_gnd_net_),
            .in3(N__26764),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__30100),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_11_13_3  (
            .in0(N__26734),
            .in1(N__26706),
            .in2(_gnd_net_),
            .in3(N__30327),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__30100),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_11_13_4  (
            .in0(N__30326),
            .in1(N__26656),
            .in2(_gnd_net_),
            .in3(N__26629),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__30100),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_11_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_11_14_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_11_14_0  (
            .in0(N__33853),
            .in1(N__33873),
            .in2(N__27169),
            .in3(N__27241),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_11_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_11_14_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_11_14_1  (
            .in0(N__27240),
            .in1(N__33852),
            .in2(N__33877),
            .in3(N__27165),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_11_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_11_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_11_14_2  (
            .in0(N__27286),
            .in1(N__27256),
            .in2(_gnd_net_),
            .in3(N__30322),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49910),
            .ce(N__30098),
            .sr(N__49459));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_11_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_11_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_11_14_3  (
            .in0(N__30321),
            .in1(N__27232),
            .in2(_gnd_net_),
            .in3(N__27207),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49910),
            .ce(N__30098),
            .sr(N__49459));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_11_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_11_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_11_14_4  (
            .in0(N__27117),
            .in1(N__27153),
            .in2(_gnd_net_),
            .in3(N__30320),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_11_15_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_11_15_0  (
            .in0(N__33805),
            .in1(N__33828),
            .in2(N__27019),
            .in3(N__27097),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_11_15_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_11_15_1  (
            .in0(N__27096),
            .in1(N__33804),
            .in2(N__33832),
            .in3(N__27015),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_11_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_11_15_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_11_15_3  (
            .in0(N__27085),
            .in1(N__27058),
            .in2(_gnd_net_),
            .in3(N__30562),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(N__30096),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_11_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_11_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_11_15_4  (
            .in0(N__30561),
            .in1(N__27006),
            .in2(_gnd_net_),
            .in3(N__26971),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(N__30096),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_15_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_15_5  (
            .in0(N__30021),
            .in1(N__30006),
            .in2(N__34102),
            .in3(N__34129),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_16_0  (
            .in0(N__31162),
            .in1(N__35542),
            .in2(N__35147),
            .in3(N__31120),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_11_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_11_16_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_11_16_1  (
            .in0(N__35539),
            .in1(N__35013),
            .in2(N__31873),
            .in3(N__31894),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_11_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_11_16_2  (
            .in0(N__32775),
            .in1(N__27478),
            .in2(_gnd_net_),
            .in3(N__28241),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_11_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_11_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_11_16_3  (
            .in0(N__35540),
            .in1(N__35014),
            .in2(N__31729),
            .in3(N__31683),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_11_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_11_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_11_16_4  (
            .in0(N__32776),
            .in1(N__31778),
            .in2(_gnd_net_),
            .in3(N__31818),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_11_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_11_16_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_11_16_5  (
            .in0(N__35544),
            .in1(N__35016),
            .in2(N__27415),
            .in3(N__28522),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_16_6  (
            .in0(N__31084),
            .in1(N__35541),
            .in2(N__35146),
            .in3(N__30912),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_16_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_16_7  (
            .in0(N__35543),
            .in1(N__35015),
            .in2(N__32395),
            .in3(N__32424),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_17_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_17_0  (
            .in0(N__28300),
            .in1(N__35453),
            .in2(N__35072),
            .in3(N__27340),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_17_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_17_1  (
            .in0(N__35450),
            .in1(N__34901),
            .in2(N__30865),
            .in3(N__30814),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_17_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_17_2  (
            .in0(N__34895),
            .in1(N__35452),
            .in2(N__31603),
            .in3(N__31641),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_11_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_11_17_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_11_17_3  (
            .in0(N__35451),
            .in1(N__34902),
            .in2(N__31369),
            .in3(N__31400),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_17_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_17_4  (
            .in0(N__34896),
            .in1(N__35454),
            .in2(N__35290),
            .in3(N__34645),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_5  (
            .in0(N__35455),
            .in1(N__34900),
            .in2(N__32074),
            .in3(N__32037),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_17_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_17_6  (
            .in0(N__34893),
            .in1(N__35456),
            .in2(N__28819),
            .in3(N__28864),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_17_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_17_7  (
            .in0(N__35449),
            .in1(N__34894),
            .in2(N__32155),
            .in3(N__32112),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__27525),
            .in2(N__27508),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__32834),
            .in2(N__32803),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__34921),
            .in2(N__31417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__30937),
            .in2(N__35108),
            .in3(N__27706),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__34925),
            .in2(N__31174),
            .in3(N__27691),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__27688),
            .in2(N__35109),
            .in3(N__27670),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__34929),
            .in2(N__31924),
            .in3(N__27655),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_11_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_11_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__31315),
            .in2(N__35110),
            .in3(N__27637),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_11_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__34933),
            .in2(N__31906),
            .in3(N__27619),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_11_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__32332),
            .in2(N__35111),
            .in3(N__27598),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_11_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__34937),
            .in2(N__32083),
            .in3(N__27586),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_11_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__32440),
            .in2(N__35112),
            .in3(N__27853),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_11_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__34941),
            .in2(N__31654),
            .in3(N__27835),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_11_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__27832),
            .in2(N__35113),
            .in3(N__27814),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_11_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_11_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__34945),
            .in2(N__30877),
            .in3(N__27799),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_11_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_11_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__31090),
            .in2(N__35114),
            .in3(N__27781),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_11_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_11_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__35115),
            .in2(N__30781),
            .in3(N__27763),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_11_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_11_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__31321),
            .in2(N__35222),
            .in3(N__27742),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_11_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_11_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__35119),
            .in2(N__30709),
            .in3(N__27724),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_11_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_11_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__31570),
            .in2(N__35223),
            .in3(N__28015),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__35123),
            .in2(N__28012),
            .in3(N__27991),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__32353),
            .in2(N__35224),
            .in3(N__27976),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__35127),
            .in2(N__27973),
            .in3(N__27946),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(N__34609),
            .in2(N__35225),
            .in3(N__27931),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__35131),
            .in2(N__31999),
            .in3(N__27916),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__35140),
            .in2(N__31495),
            .in3(N__27901),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__35132),
            .in2(N__27898),
            .in3(N__27871),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__35141),
            .in2(N__28789),
            .in3(N__28126),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__35133),
            .in2(N__31237),
            .in3(N__28111),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__35142),
            .in2(N__28714),
            .in3(N__28093),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__35134),
            .in2(N__32512),
            .in3(N__28075),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_21_7  (
            .in0(N__35135),
            .in1(N__35601),
            .in2(_gnd_net_),
            .in3(N__28072),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__32851),
            .in2(N__32247),
            .in3(N__32237),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__28057),
            .in2(_gnd_net_),
            .in3(N__28051),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__28048),
            .in2(_gnd_net_),
            .in3(N__28042),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__28039),
            .in2(_gnd_net_),
            .in3(N__28033),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__28261),
            .in2(_gnd_net_),
            .in3(N__28219),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__28216),
            .in2(_gnd_net_),
            .in3(N__28210),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__28207),
            .in2(_gnd_net_),
            .in3(N__28198),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__28195),
            .in2(_gnd_net_),
            .in3(N__28186),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__28183),
            .in2(_gnd_net_),
            .in3(N__28174),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__28171),
            .in2(_gnd_net_),
            .in3(N__28165),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__28162),
            .in2(_gnd_net_),
            .in3(N__28150),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__28147),
            .in2(_gnd_net_),
            .in3(N__28141),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__28393),
            .in2(_gnd_net_),
            .in3(N__28360),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__31042),
            .in2(_gnd_net_),
            .in3(N__28357),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__28354),
            .in2(_gnd_net_),
            .in3(N__28348),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(N__28345),
            .in2(_gnd_net_),
            .in3(N__28339),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__28336),
            .in2(_gnd_net_),
            .in3(N__28327),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__28324),
            .in2(_gnd_net_),
            .in3(N__28318),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__28315),
            .in2(_gnd_net_),
            .in3(N__28309),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__28306),
            .in2(_gnd_net_),
            .in3(N__28273),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__28270),
            .in2(_gnd_net_),
            .in3(N__28264),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__28528),
            .in2(_gnd_net_),
            .in3(N__28495),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__28492),
            .in2(_gnd_net_),
            .in3(N__28486),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__28483),
            .in2(_gnd_net_),
            .in3(N__28477),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__28474),
            .in2(_gnd_net_),
            .in3(N__28468),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_25_1  (
            .in0(_gnd_net_),
            .in1(N__28465),
            .in2(_gnd_net_),
            .in3(N__28429),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(N__28426),
            .in2(_gnd_net_),
            .in3(N__28414),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(N__28411),
            .in2(_gnd_net_),
            .in3(N__28405),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__28402),
            .in2(_gnd_net_),
            .in3(N__28396),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28867),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_25_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_25_6  (
            .in0(N__35610),
            .in1(N__35244),
            .in2(N__28863),
            .in3(N__28808),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_25_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_25_7  (
            .in0(N__35245),
            .in1(N__35611),
            .in2(N__28777),
            .in3(N__28733),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_11_27_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_11_27_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_11_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_11_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42013),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49867),
            .ce(),
            .sr(N__49523));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28687),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_12_6_0  (
            .in0(N__28667),
            .in1(N__28651),
            .in2(_gnd_net_),
            .in3(N__30424),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49967),
            .ce(N__30106),
            .sr(N__49392));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_7_3 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_12_7_3  (
            .in0(N__39996),
            .in1(N__28609),
            .in2(N__28585),
            .in3(N__28555),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49958),
            .ce(),
            .sr(N__49398));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_12_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_12_8_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_12_8_0  (
            .in0(N__43448),
            .in1(N__43415),
            .in2(N__48392),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_12_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_12_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_12_8_1  (
            .in0(N__43799),
            .in1(N__43779),
            .in2(_gnd_net_),
            .in3(N__48362),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_12_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_12_8_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_12_8_2  (
            .in0(N__44000),
            .in1(N__44024),
            .in2(N__48391),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_12_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_12_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_12_8_4  (
            .in0(N__29537),
            .in1(N__29517),
            .in2(_gnd_net_),
            .in3(N__30498),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_12_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_12_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_12_9_0  (
            .in0(N__28907),
            .in1(N__28878),
            .in2(_gnd_net_),
            .in3(N__30490),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_9_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_12_9_1  (
            .in0(N__30491),
            .in1(_gnd_net_),
            .in2(N__29302),
            .in3(N__28908),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49941),
            .ce(N__29253),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_12_9_2  (
            .in0(N__29395),
            .in1(N__29410),
            .in2(_gnd_net_),
            .in3(N__30492),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49941),
            .ce(N__29253),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_12_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_12_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_12_9_5  (
            .in0(N__48358),
            .in1(N__44159),
            .in2(_gnd_net_),
            .in3(N__44135),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_9_7  (
            .in0(N__28999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48570),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_12_10_3  (
            .in0(N__28951),
            .in1(N__28924),
            .in2(_gnd_net_),
            .in3(N__30555),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(N__30105),
            .sr(N__49417));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_12_10_5  (
            .in0(N__28909),
            .in1(N__28879),
            .in2(_gnd_net_),
            .in3(N__30556),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(N__30105),
            .sr(N__49417));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_12_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_12_10_6  (
            .in0(N__30554),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(N__29518),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(N__30105),
            .sr(N__49417));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_11_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_11_0  (
            .in0(N__33561),
            .in1(N__29419),
            .in2(N__29476),
            .in3(N__33903),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_11_1  (
            .in0(N__29418),
            .in1(N__33562),
            .in2(N__33904),
            .in3(N__29475),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_12_11_2  (
            .in0(N__29464),
            .in1(N__29434),
            .in2(_gnd_net_),
            .in3(N__30435),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(N__30104),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_12_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_12_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_12_11_4  (
            .in0(N__29393),
            .in1(N__29406),
            .in2(_gnd_net_),
            .in3(N__30433),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_11_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_12_11_5  (
            .in0(N__30434),
            .in1(N__29394),
            .in2(N__29365),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(N__30104),
            .sr(N__49425));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_12_11_6  (
            .in0(N__29362),
            .in1(N__29332),
            .in2(_gnd_net_),
            .in3(N__30436),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(N__30104),
            .sr(N__49425));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__29308),
            .in2(N__29320),
            .in3(N__41538),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__29674),
            .in2(N__29668),
            .in3(N__33378),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__29659),
            .in2(N__29647),
            .in3(N__33360),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__29638),
            .in2(N__29629),
            .in3(N__33540),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__29620),
            .in2(N__29614),
            .in3(N__33526),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__29593),
            .in2(N__29602),
            .in3(N__33507),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__29578),
            .in2(N__29587),
            .in3(N__33492),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__29563),
            .in2(N__29572),
            .in3(N__33477),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__29557),
            .in2(N__29548),
            .in3(N__33463),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_13_1  (
            .in0(N__33445),
            .in1(N__29809),
            .in2(N__29821),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__29791),
            .in2(N__29803),
            .in3(N__33426),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__29785),
            .in2(N__29776),
            .in3(N__33411),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(N__29752),
            .in3(N__33708),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__29743),
            .in2(N__29734),
            .in3(N__33693),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__29725),
            .in2(N__29716),
            .in3(N__33678),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__29707),
            .in2(N__29701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__29692),
            .in2(N__29686),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__29896),
            .in2(N__29887),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__29875),
            .in2(N__29866),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__29854),
            .in2(N__29848),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__30682),
            .in2(N__29830),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__30067),
            .in2(N__30034),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_12_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_12_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__29839),
            .in2(N__29992),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29833),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_12_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_12_15_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_12_15_0  (
            .in0(N__33783),
            .in1(N__30696),
            .in2(N__33766),
            .in3(N__30628),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_15_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_15_1  (
            .in0(N__30627),
            .in1(N__33761),
            .in2(N__30700),
            .in3(N__33782),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_12_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_12_15_2  (
            .in0(N__30676),
            .in1(N__30646),
            .in2(_gnd_net_),
            .in3(N__30559),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(N__30099),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_12_15_4  (
            .in0(N__30619),
            .in1(N__30580),
            .in2(_gnd_net_),
            .in3(N__30560),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(N__30099),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_15_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_15_5  (
            .in0(N__30042),
            .in1(N__33722),
            .in2(N__30061),
            .in3(N__33743),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_15_6 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_15_6  (
            .in0(N__33723),
            .in1(N__30057),
            .in2(N__33745),
            .in3(N__30043),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_16_1 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_16_1  (
            .in0(N__30025),
            .in1(N__34097),
            .in2(N__30007),
            .in3(N__34127),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29979),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49472));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29953),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49472));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_12_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_12_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_12_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29925),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49472));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31030),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49472));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_12_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_12_18_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_12_18_4  (
            .in0(N__35186),
            .in1(N__35423),
            .in2(N__30987),
            .in3(N__30957),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32188),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__32878),
            .sr(N__49479));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_12_18_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_12_18_6  (
            .in0(N__35187),
            .in1(N__35424),
            .in2(N__30988),
            .in3(N__30958),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_7  (
            .in0(N__35422),
            .in1(N__35188),
            .in2(N__31482),
            .in3(N__31441),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_12_19_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_12_19_0  (
            .in0(N__35426),
            .in1(N__35227),
            .in2(N__30913),
            .in3(N__31080),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_12_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_12_19_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_12_19_1  (
            .in0(N__35228),
            .in1(N__35427),
            .in2(N__30864),
            .in3(N__30813),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_12_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_12_19_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_12_19_2  (
            .in0(N__35429),
            .in1(N__35226),
            .in2(N__30772),
            .in3(N__30733),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_12_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_12_19_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_12_19_4  (
            .in0(N__35430),
            .in1(N__35229),
            .in2(N__31564),
            .in3(N__31528),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_19_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_19_6  (
            .in0(N__35425),
            .in1(N__35231),
            .in2(N__31483),
            .in3(N__31437),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_12_19_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_12_19_7  (
            .in0(N__35230),
            .in1(N__35428),
            .in2(N__31405),
            .in3(N__31365),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_20_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_20_0  (
            .in0(N__35497),
            .in1(N__35175),
            .in2(N__31782),
            .in3(N__31819),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_12_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_12_20_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_12_20_1  (
            .in0(N__31306),
            .in1(N__35501),
            .in2(N__35234),
            .in3(N__31270),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_12_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_12_20_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_12_20_3  (
            .in0(N__31228),
            .in1(N__35496),
            .in2(N__35233),
            .in3(N__31201),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_20_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_20_4  (
            .in0(N__35499),
            .in1(N__35176),
            .in2(N__31161),
            .in3(N__31119),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31072),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_12_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_12_20_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_12_20_6  (
            .in0(N__35498),
            .in1(N__35171),
            .in2(N__32151),
            .in3(N__32111),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_12_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_12_20_7 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_12_20_7  (
            .in0(N__35177),
            .in1(N__32067),
            .in2(N__32041),
            .in3(N__35500),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_21_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_21_0  (
            .in0(N__35562),
            .in1(N__35215),
            .in2(N__31990),
            .in3(N__31960),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_21_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_21_1  (
            .in0(N__35218),
            .in1(N__35564),
            .in2(N__31872),
            .in3(N__31887),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_12_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_12_21_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_12_21_2  (
            .in0(N__31886),
            .in1(N__32704),
            .in2(_gnd_net_),
            .in3(N__31865),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_12_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_12_21_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_12_21_3  (
            .in0(N__35216),
            .in1(N__35563),
            .in2(N__31814),
            .in3(N__31786),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_21_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_21_4  (
            .in0(N__35566),
            .in1(N__35219),
            .in2(N__31722),
            .in3(N__31682),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_12_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_12_21_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_12_21_5  (
            .in0(N__35221),
            .in1(N__35567),
            .in2(N__31642),
            .in3(N__31598),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_12_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_12_21_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_12_21_6  (
            .in0(N__35565),
            .in1(N__32494),
            .in2(N__32470),
            .in3(N__35217),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_12_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_12_21_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_12_21_7  (
            .in0(N__35220),
            .in1(N__35568),
            .in2(N__32428),
            .in3(N__32391),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_22_0 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_22_0  (
            .in0(N__32274),
            .in1(N__35569),
            .in2(N__32305),
            .in3(N__35164),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_12_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_12_22_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_12_22_1  (
            .in0(N__35570),
            .in1(N__32304),
            .in2(N__35232),
            .in3(N__32275),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_12_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_12_22_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__35571),
            .in2(_gnd_net_),
            .in3(N__35163),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_12_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_12_22_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_12_22_3  (
            .in0(N__32300),
            .in1(N__32683),
            .in2(_gnd_net_),
            .in3(N__32273),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32939),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_12_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_12_22_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_12_22_5  (
            .in0(N__32940),
            .in1(_gnd_net_),
            .in2(N__32218),
            .in3(N__32682),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_12_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_12_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_12_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32184),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__32875),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32977),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__32875),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_23_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_23_0  (
            .in0(N__35536),
            .in1(N__32643),
            .in2(N__32839),
            .in3(N__32631),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32905),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49873),
            .ce(N__32874),
            .sr(N__49502));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32629),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_23_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_23_3  (
            .in0(N__32632),
            .in1(N__35537),
            .in2(N__32647),
            .in3(N__32838),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_23_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_23_4  (
            .in0(N__32684),
            .in1(N__32642),
            .in2(_gnd_net_),
            .in3(N__32630),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_12_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_12_23_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_12_23_6  (
            .in0(N__35538),
            .in1(N__35236),
            .in2(N__32599),
            .in3(N__32534),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_12_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_12_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__34527),
            .in2(_gnd_net_),
            .in3(N__34593),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_12_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_12_24_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_12_24_1  (
            .in0(N__34468),
            .in1(N__34495),
            .in2(N__32497),
            .in3(N__34564),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_12_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_12_25_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_12_25_3  (
            .in0(N__35706),
            .in1(N__35733),
            .in2(_gnd_net_),
            .in3(N__35759),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_12_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_12_25_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_12_25_4  (
            .in0(N__35787),
            .in1(N__33007),
            .in2(N__33001),
            .in3(N__34437),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_12_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_12_26_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_12_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_12_26_0  (
            .in0(N__33071),
            .in1(N__34592),
            .in2(_gnd_net_),
            .in3(N__32998),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_26_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_1_LC_12_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_12_26_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_12_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_12_26_1  (
            .in0(N__33067),
            .in1(N__34556),
            .in2(_gnd_net_),
            .in3(N__32995),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_2_LC_12_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_12_26_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_12_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_12_26_2  (
            .in0(N__33072),
            .in1(N__34526),
            .in2(_gnd_net_),
            .in3(N__32992),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_3_LC_12_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_12_26_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_12_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_12_26_3  (
            .in0(N__33068),
            .in1(N__34493),
            .in2(_gnd_net_),
            .in3(N__32989),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_4_LC_12_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_12_26_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_12_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_12_26_4  (
            .in0(N__33073),
            .in1(N__34466),
            .in2(_gnd_net_),
            .in3(N__32986),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_5_LC_12_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_12_26_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_12_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_12_26_5  (
            .in0(N__33069),
            .in1(N__34436),
            .in2(_gnd_net_),
            .in3(N__32983),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_6_LC_12_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_12_26_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_12_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_12_26_6  (
            .in0(N__33074),
            .in1(N__35786),
            .in2(_gnd_net_),
            .in3(N__32980),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_7_LC_12_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_12_26_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_12_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_12_26_7  (
            .in0(N__33070),
            .in1(N__35760),
            .in2(_gnd_net_),
            .in3(N__33082),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49517));
    defparam \pwm_generator_inst.counter_8_LC_12_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_12_27_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_12_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_12_27_0  (
            .in0(N__33076),
            .in1(N__35732),
            .in2(_gnd_net_),
            .in3(N__33079),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__49865),
            .ce(),
            .sr(N__49521));
    defparam \pwm_generator_inst.counter_9_LC_12_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_12_27_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_12_27_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_12_27_1  (
            .in0(N__35705),
            .in1(N__33075),
            .in2(_gnd_net_),
            .in3(N__33034),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49865),
            .ce(),
            .sr(N__49521));
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_6.C_ON=1'b0;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_6 (
            .in0(N__49552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_red_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_6_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__36009),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49978),
            .ce(N__36462),
            .sr(N__49385));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_6_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__35988),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49978),
            .ce(N__36462),
            .sr(N__49385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_7_0  (
            .in0(N__33320),
            .in1(N__36005),
            .in2(_gnd_net_),
            .in3(N__33016),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_7_1  (
            .in0(N__33315),
            .in1(N__35984),
            .in2(_gnd_net_),
            .in3(N__33013),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_7_2  (
            .in0(N__33321),
            .in1(N__35961),
            .in2(_gnd_net_),
            .in3(N__33010),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_7_3  (
            .in0(N__33316),
            .in1(N__35937),
            .in2(_gnd_net_),
            .in3(N__33109),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_7_4  (
            .in0(N__33322),
            .in1(N__35913),
            .in2(_gnd_net_),
            .in3(N__33106),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_7_5  (
            .in0(N__33317),
            .in1(N__35889),
            .in2(_gnd_net_),
            .in3(N__33103),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_7_6  (
            .in0(N__33319),
            .in1(N__35865),
            .in2(_gnd_net_),
            .in3(N__33100),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_7_7  (
            .in0(N__33318),
            .in1(N__35841),
            .in2(_gnd_net_),
            .in3(N__33097),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49969),
            .ce(N__33187),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_8_0  (
            .in0(N__33311),
            .in1(N__36198),
            .in2(_gnd_net_),
            .in3(N__33094),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_8_1  (
            .in0(N__33296),
            .in1(N__36174),
            .in2(_gnd_net_),
            .in3(N__33091),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_8_2  (
            .in0(N__33308),
            .in1(N__36150),
            .in2(_gnd_net_),
            .in3(N__33088),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_8_3  (
            .in0(N__33293),
            .in1(N__36126),
            .in2(_gnd_net_),
            .in3(N__33085),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_8_4  (
            .in0(N__33309),
            .in1(N__36102),
            .in2(_gnd_net_),
            .in3(N__33136),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_8_5  (
            .in0(N__33294),
            .in1(N__36078),
            .in2(_gnd_net_),
            .in3(N__33133),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_8_6  (
            .in0(N__33310),
            .in1(N__36054),
            .in2(_gnd_net_),
            .in3(N__33130),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_8_7  (
            .in0(N__33295),
            .in1(N__36030),
            .in2(_gnd_net_),
            .in3(N__33127),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49960),
            .ce(N__33182),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_9_0  (
            .in0(N__33297),
            .in1(N__36387),
            .in2(_gnd_net_),
            .in3(N__33124),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_9_1  (
            .in0(N__33301),
            .in1(N__36363),
            .in2(_gnd_net_),
            .in3(N__33121),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_9_2  (
            .in0(N__33298),
            .in1(N__36343),
            .in2(_gnd_net_),
            .in3(N__33118),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_9_3  (
            .in0(N__33302),
            .in1(N__36321),
            .in2(_gnd_net_),
            .in3(N__33115),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_9_4  (
            .in0(N__33299),
            .in1(N__36299),
            .in2(_gnd_net_),
            .in3(N__33112),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_9_5  (
            .in0(N__33303),
            .in1(N__36273),
            .in2(_gnd_net_),
            .in3(N__33346),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_9_6  (
            .in0(N__33300),
            .in1(N__36249),
            .in2(_gnd_net_),
            .in3(N__33343),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_9_7  (
            .in0(N__33304),
            .in1(N__36225),
            .in2(_gnd_net_),
            .in3(N__33340),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49951),
            .ce(N__33181),
            .sr(N__49405));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_10_0  (
            .in0(N__33312),
            .in1(N__36582),
            .in2(_gnd_net_),
            .in3(N__33337),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_10_1  (
            .in0(N__33305),
            .in1(N__36558),
            .in2(_gnd_net_),
            .in3(N__33334),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_10_2  (
            .in0(N__33313),
            .in1(N__36522),
            .in2(_gnd_net_),
            .in3(N__33331),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_10_3  (
            .in0(N__33306),
            .in1(N__36486),
            .in2(_gnd_net_),
            .in3(N__33328),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_10_4  (
            .in0(N__33314),
            .in1(N__36538),
            .in2(_gnd_net_),
            .in3(N__33325),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_10_5  (
            .in0(N__33307),
            .in1(N__36502),
            .in2(_gnd_net_),
            .in3(N__33190),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(N__33186),
            .sr(N__49411));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_13_11_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_13_11_0  (
            .in0(N__33397),
            .in1(N__39829),
            .in2(N__39805),
            .in3(N__33388),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_13_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_13_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_13_11_2  (
            .in0(N__41518),
            .in1(N__41489),
            .in2(_gnd_net_),
            .in3(N__48398),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(N__45840),
            .sr(N__49418));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_13_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_13_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_13_11_3  (
            .in0(N__48397),
            .in1(N__41431),
            .in2(_gnd_net_),
            .in3(N__41407),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(N__45840),
            .sr(N__49418));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_13_11_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_13_11_4  (
            .in0(N__33396),
            .in1(N__39828),
            .in2(N__39804),
            .in3(N__33387),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_13_11_6  (
            .in0(N__47524),
            .in1(N__47500),
            .in2(_gnd_net_),
            .in3(N__48399),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(N__45840),
            .sr(N__49418));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_7 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_7  (
            .in0(N__36645),
            .in1(N__39687),
            .in2(N__39724),
            .in3(N__36633),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_13_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_13_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__41539),
            .in2(N__36622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_13_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_13_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_13_12_1  (
            .in0(N__41230),
            .in1(N__33379),
            .in2(_gnd_net_),
            .in3(N__33367),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_13_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_13_12_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_13_12_2  (
            .in0(N__41260),
            .in1(N__36607),
            .in2(N__33364),
            .in3(N__33349),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_13_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_13_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_13_12_3  (
            .in0(N__41231),
            .in1(N__33541),
            .in2(_gnd_net_),
            .in3(N__33529),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_13_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_13_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_13_12_4  (
            .in0(N__41261),
            .in1(N__33525),
            .in2(_gnd_net_),
            .in3(N__33511),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_13_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_13_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_13_12_5  (
            .in0(N__41232),
            .in1(N__33508),
            .in2(_gnd_net_),
            .in3(N__33496),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_13_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_13_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_13_12_6  (
            .in0(N__41262),
            .in1(N__33493),
            .in2(_gnd_net_),
            .in3(N__33481),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_13_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_13_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_13_12_7  (
            .in0(N__41233),
            .in1(N__33478),
            .in2(_gnd_net_),
            .in3(N__33466),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_13_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_13_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_13_13_0  (
            .in0(N__41255),
            .in1(N__33462),
            .in2(_gnd_net_),
            .in3(N__33448),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_13_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_13_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_13_13_1  (
            .in0(N__41256),
            .in1(N__33444),
            .in2(_gnd_net_),
            .in3(N__33430),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_13_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_13_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_13_13_2  (
            .in0(N__41252),
            .in1(N__33427),
            .in2(_gnd_net_),
            .in3(N__33415),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_13_3  (
            .in0(N__41257),
            .in1(N__33412),
            .in2(_gnd_net_),
            .in3(N__33400),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_13_4  (
            .in0(N__41253),
            .in1(N__33709),
            .in2(_gnd_net_),
            .in3(N__33697),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_13_5  (
            .in0(N__41258),
            .in1(N__33694),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_13_6  (
            .in0(N__41254),
            .in1(N__33679),
            .in2(_gnd_net_),
            .in3(N__33667),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_13_7  (
            .in0(N__41259),
            .in1(N__33657),
            .in2(_gnd_net_),
            .in3(N__33643),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49915),
            .ce(),
            .sr(N__49433));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_14_0  (
            .in0(N__41240),
            .in1(N__33630),
            .in2(_gnd_net_),
            .in3(N__33616),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_14_1  (
            .in0(N__41244),
            .in1(N__33603),
            .in2(_gnd_net_),
            .in3(N__33589),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_14_2  (
            .in0(N__41241),
            .in1(N__33579),
            .in2(_gnd_net_),
            .in3(N__33565),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_13_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_13_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_13_14_3  (
            .in0(N__41245),
            .in1(N__33560),
            .in2(_gnd_net_),
            .in3(N__33544),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_13_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_13_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_13_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_13_14_4  (
            .in0(N__41242),
            .in1(N__33894),
            .in2(_gnd_net_),
            .in3(N__33880),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_13_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_13_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_13_14_5  (
            .in0(N__41246),
            .in1(N__33872),
            .in2(_gnd_net_),
            .in3(N__33856),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_13_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_13_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_13_14_6  (
            .in0(N__41243),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__33835),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_13_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_13_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_13_14_7  (
            .in0(N__41247),
            .in1(N__33822),
            .in2(_gnd_net_),
            .in3(N__33808),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49911),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_13_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_13_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_13_15_0  (
            .in0(N__41248),
            .in1(N__33803),
            .in2(_gnd_net_),
            .in3(N__33787),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_13_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_13_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_13_15_1  (
            .in0(N__41237),
            .in1(N__33784),
            .in2(_gnd_net_),
            .in3(N__33769),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_13_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_13_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_13_15_2  (
            .in0(N__41249),
            .in1(N__33765),
            .in2(_gnd_net_),
            .in3(N__33748),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_13_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_13_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_13_15_3  (
            .in0(N__41238),
            .in1(N__33744),
            .in2(_gnd_net_),
            .in3(N__33727),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_13_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_13_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_13_15_4  (
            .in0(N__41250),
            .in1(N__33724),
            .in2(_gnd_net_),
            .in3(N__34132),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_13_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_13_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_13_15_5  (
            .in0(N__41239),
            .in1(N__34128),
            .in2(_gnd_net_),
            .in3(N__34108),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_13_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_13_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_13_15_6  (
            .in0(N__41251),
            .in1(N__34098),
            .in2(_gnd_net_),
            .in3(N__34105),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49905),
            .ce(),
            .sr(N__49451));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34078),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49900),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34048),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49900),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49900),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_13_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_13_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33994),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49900),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33964),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49896),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33936),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49896),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34411),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49896),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34384),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49896),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34353),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49473));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34329),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49473));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_13_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34300),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49473));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34272),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49885),
            .ce(),
            .sr(N__49480));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34242),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49885),
            .ce(),
            .sr(N__49480));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34209),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49885),
            .ce(),
            .sr(N__49480));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34176),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49885),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst1.S2_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.S2_LC_13_20_0  (
            .in0(N__41626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49880),
            .ce(),
            .sr(N__49485));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35643),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49880),
            .ce(),
            .sr(N__49485));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_22_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_22_6  (
            .in0(N__35572),
            .in1(N__35279),
            .in2(N__35235),
            .in3(N__34638),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__34570),
            .in2(N__38857),
            .in3(N__34597),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__38557),
            .in2(N__34540),
            .in3(N__34563),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__38887),
            .in2(N__34504),
            .in3(N__34531),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__34474),
            .in2(N__38572),
            .in3(N__34494),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4  (
            .in0(N__34467),
            .in1(N__38587),
            .in2(N__34447),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5  (
            .in0(N__34438),
            .in1(N__34417),
            .in2(N__38542),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6  (
            .in0(N__35788),
            .in1(N__35767),
            .in2(N__38602),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7  (
            .in0(N__35761),
            .in1(N__35740),
            .in2(N__38872),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__35713),
            .in2(N__38839),
            .in3(N__35734),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__35683),
            .in2(N__35800),
            .in3(N__35707),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35677),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(),
            .sr(N__49508));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__38830),
            .in2(N__44989),
            .in3(N__44976),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__44866),
            .in2(_gnd_net_),
            .in3(N__35650),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__38818),
            .in2(_gnd_net_),
            .in3(N__35647),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__38824),
            .in2(_gnd_net_),
            .in3(N__35824),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__38812),
            .in2(_gnd_net_),
            .in3(N__35821),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__42169),
            .in2(_gnd_net_),
            .in3(N__35818),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__43219),
            .in2(_gnd_net_),
            .in3(N__35815),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__38926),
            .in2(_gnd_net_),
            .in3(N__35812),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__43231),
            .in2(_gnd_net_),
            .in3(N__35809),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_13_27_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_27_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_27_1  (
            .in0(N__45166),
            .in1(N__40396),
            .in2(N__44992),
            .in3(N__35806),
            .lcout(),
            .ltout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_13_27_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_13_27_2 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_13_27_2  (
            .in0(N__49051),
            .in1(N__47848),
            .in2(N__35803),
            .in3(N__42312),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_14_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_14_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_14_5_3  (
            .in0(N__44091),
            .in1(N__44069),
            .in2(_gnd_net_),
            .in3(N__48329),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_14_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_14_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_14_6_6  (
            .in0(N__45536),
            .in1(N__45509),
            .in2(_gnd_net_),
            .in3(N__48348),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__35960),
            .in2(N__36010),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__35936),
            .in2(N__35989),
            .in3(N__35968),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__35912),
            .in2(N__35965),
            .in3(N__35944),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__35888),
            .in2(N__35941),
            .in3(N__35920),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__35864),
            .in2(N__35917),
            .in3(N__35896),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__35840),
            .in2(N__35893),
            .in3(N__35872),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__36197),
            .in2(N__35869),
            .in3(N__35848),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__36173),
            .in2(N__35845),
            .in3(N__36205),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49979),
            .ce(N__36463),
            .sr(N__49386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__36149),
            .in2(N__36202),
            .in3(N__36181),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__36125),
            .in2(N__36178),
            .in3(N__36157),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__36101),
            .in2(N__36154),
            .in3(N__36133),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__36077),
            .in2(N__36130),
            .in3(N__36109),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__36053),
            .in2(N__36106),
            .in3(N__36085),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__36029),
            .in2(N__36082),
            .in3(N__36061),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__36386),
            .in2(N__36058),
            .in3(N__36037),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__36362),
            .in2(N__36034),
            .in3(N__36013),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49970),
            .ce(N__36461),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__36341),
            .in2(N__36391),
            .in3(N__36370),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__36320),
            .in2(N__36367),
            .in3(N__36346),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__36342),
            .in2(N__36300),
            .in3(N__36328),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__36272),
            .in2(N__36325),
            .in3(N__36304),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__36248),
            .in2(N__36301),
            .in3(N__36280),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__36224),
            .in2(N__36277),
            .in3(N__36256),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__36581),
            .in2(N__36253),
            .in3(N__36232),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__36557),
            .in2(N__36229),
            .in3(N__36208),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49961),
            .ce(N__36447),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__36521),
            .in2(N__36586),
            .in3(N__36565),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49952),
            .ce(N__36460),
            .sr(N__49406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__36485),
            .in2(N__36562),
            .in3(N__36541),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49952),
            .ce(N__36460),
            .sr(N__49406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__36537),
            .in2(N__36526),
            .in3(N__36505),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49952),
            .ce(N__36460),
            .sr(N__49406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__36501),
            .in2(N__36490),
            .in3(N__36469),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49952),
            .ce(N__36460),
            .sr(N__49406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36466),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(N__36460),
            .sr(N__49406));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_14_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_14_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_14_11_0  (
            .in0(N__39748),
            .in1(N__39771),
            .in2(N__36403),
            .in3(N__36655),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_14_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_14_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_14_11_1  (
            .in0(N__36654),
            .in1(N__39747),
            .in2(N__39775),
            .in3(N__36399),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_14_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_14_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_14_11_2  (
            .in0(N__41879),
            .in1(N__48393),
            .in2(_gnd_net_),
            .in3(N__41898),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_14_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_14_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_14_11_3  (
            .in0(N__48395),
            .in1(_gnd_net_),
            .in2(N__36406),
            .in3(N__41880),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(N__45844),
            .sr(N__49412));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_14_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_14_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_14_11_5  (
            .in0(N__48394),
            .in1(N__46168),
            .in2(_gnd_net_),
            .in3(N__46146),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(N__45844),
            .sr(N__49412));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_14_11_6  (
            .in0(N__48613),
            .in1(N__48649),
            .in2(_gnd_net_),
            .in3(N__48396),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(N__45844),
            .sr(N__49412));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_14_11_7 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_14_11_7  (
            .in0(N__36646),
            .in1(N__39723),
            .in2(N__39691),
            .in3(N__36634),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__41582),
            .in2(_gnd_net_),
            .in3(N__41553),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_14_12_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__41303),
            .in2(_gnd_net_),
            .in3(N__36771),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_14_12_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36610),
            .in3(N__41583),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_14_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_14_13_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_14_13_0  (
            .in0(N__36793),
            .in1(N__39568),
            .in2(N__36601),
            .in3(N__39585),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_14_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_14_13_3  (
            .in0(N__47632),
            .in1(N__47593),
            .in2(_gnd_net_),
            .in3(N__48383),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(N__45835),
            .sr(N__49427));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_13_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_13_4  (
            .in0(N__36792),
            .in1(N__39567),
            .in2(N__36600),
            .in3(N__39584),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_14_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_14_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_14_13_5  (
            .in0(N__47722),
            .in1(N__47689),
            .in2(_gnd_net_),
            .in3(N__48382),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(N__45835),
            .sr(N__49427));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_14_13_7  (
            .in0(N__44035),
            .in1(N__44001),
            .in2(_gnd_net_),
            .in3(N__48384),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(N__45835),
            .sr(N__49427));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_14_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_14_0  (
            .in0(N__41770),
            .in1(N__41335),
            .in2(N__39407),
            .in3(N__45828),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_14_14_3 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_14_14_3  (
            .in0(N__41295),
            .in1(N__36780),
            .in2(_gnd_net_),
            .in3(N__42147),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_LC_14_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_14_14_4 .LUT_INIT=16'b1011101000111010;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_14_14_4  (
            .in0(N__36781),
            .in1(N__41296),
            .in2(N__36784),
            .in3(N__36767),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42148),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_14_15_0 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_14_15_0  (
            .in0(N__36772),
            .in1(N__40354),
            .in2(N__41307),
            .in3(N__41578),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_14_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_14_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36741),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_14_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_14_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36715),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_14_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_14_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36685),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(),
            .sr(N__49452));
    defparam \phase_controller_inst1.state_2_LC_14_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_16_3 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_16_3  (
            .in0(N__41717),
            .in1(N__42443),
            .in2(N__40018),
            .in3(N__40035),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(),
            .sr(N__49452));
    defparam \phase_controller_inst1.start_timer_hc_LC_14_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_14_16_7 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_14_16_7  (
            .in0(N__41730),
            .in1(N__44739),
            .in2(N__37115),
            .in3(N__39658),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(),
            .sr(N__49452));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_14_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__46695),
            .in2(N__39946),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__37093),
            .in2(N__37084),
            .in3(N__37045),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__37042),
            .in2(N__37036),
            .in3(N__36985),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__36982),
            .in2(N__36976),
            .in3(N__36925),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__39952),
            .in2(N__36922),
            .in3(N__36865),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__36862),
            .in2(N__36853),
            .in3(N__36796),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__37615),
            .in2(N__37606),
            .in3(N__37555),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__37552),
            .in2(N__37546),
            .in3(N__37498),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__37495),
            .in2(N__37489),
            .in3(N__37438),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__37435),
            .in2(N__37378),
            .in3(N__37366),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__37363),
            .in2(N__37351),
            .in3(N__37306),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__37303),
            .in2(N__37294),
            .in3(N__37243),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__37240),
            .in2(N__37234),
            .in3(N__37183),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__37180),
            .in2(N__37174),
            .in3(N__37129),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__38062),
            .in2(N__38047),
            .in3(N__37999),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_14_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__37996),
            .in2(N__37990),
            .in3(N__37942),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_14_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_14_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__37939),
            .in2(N__37933),
            .in3(N__37891),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_14_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__37888),
            .in2(N__37849),
            .in3(N__37840),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_14_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__37837),
            .in2(N__37795),
            .in3(N__37783),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_14_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__37780),
            .in2(N__37774),
            .in3(N__37723),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_14_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__37720),
            .in2(N__37711),
            .in3(N__37675),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_14_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__37672),
            .in2(N__37666),
            .in3(N__37618),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_14_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__38533),
            .in2(N__38521),
            .in3(N__38473),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_14_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__38470),
            .in2(N__38461),
            .in3(N__38410),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49891),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_14_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_14_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__38407),
            .in2(N__38398),
            .in3(N__38359),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_14_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__38356),
            .in2(N__38347),
            .in3(N__38299),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_14_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__38296),
            .in2(N__38281),
            .in3(N__38233),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_14_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__38230),
            .in2(N__38191),
            .in3(N__38182),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_14_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__38179),
            .in2(N__38173),
            .in3(N__38128),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_14_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__38125),
            .in2(N__38110),
            .in3(N__38806),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_14_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_14_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_14_20_6  (
            .in0(N__38617),
            .in1(N__38801),
            .in2(_gnd_net_),
            .in3(N__38635),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_14_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_14_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_14_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38632),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(),
            .sr(N__49481));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_14_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_14_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__40383),
            .in2(_gnd_net_),
            .in3(N__40355),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_14_25_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_14_25_0 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_14_25_0  (
            .in0(N__49046),
            .in1(N__47843),
            .in2(N__38611),
            .in3(N__42310),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_14_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_14_25_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_14_25_1  (
            .in0(N__47841),
            .in1(N__38593),
            .in2(N__42359),
            .in3(N__49044),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_14_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_14_25_2 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_14_25_2  (
            .in0(N__49043),
            .in1(N__47840),
            .in2(N__38581),
            .in3(N__42305),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_14_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_14_25_3 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_14_25_3  (
            .in0(N__47838),
            .in1(N__38563),
            .in2(N__42357),
            .in3(N__49041),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_14_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_14_25_4 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_14_25_4  (
            .in0(N__49045),
            .in1(N__47842),
            .in2(N__38551),
            .in3(N__42309),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_14_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_14_25_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_14_25_5  (
            .in0(N__47839),
            .in1(N__38893),
            .in2(N__42358),
            .in3(N__49042),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_14_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_14_25_6 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_14_25_6  (
            .in0(N__49047),
            .in1(N__47844),
            .in2(N__38881),
            .in3(N__42311),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_26_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_26_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_26_5  (
            .in0(N__47818),
            .in1(N__38863),
            .in2(N__42356),
            .in3(N__49016),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_14_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_14_26_6 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_14_26_6  (
            .in0(N__49017),
            .in1(N__47819),
            .in2(N__42360),
            .in3(N__38845),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_14_27_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_14_27_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_14_27_0  (
            .in0(N__46678),
            .in1(N__46654),
            .in2(N__44990),
            .in3(N__45004),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_14_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_14_27_1 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_14_27_1  (
            .in0(N__44984),
            .in1(N__45316),
            .in2(N__42913),
            .in3(N__45340),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_14_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_14_27_3 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_14_27_3  (
            .in0(N__44983),
            .in1(N__44824),
            .in2(N__44851),
            .in3(N__42193),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_14_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_14_27_4 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_14_27_4  (
            .in0(N__45304),
            .in1(N__45280),
            .in2(N__44991),
            .in3(N__42160),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(N__40800),
            .in2(_gnd_net_),
            .in3(N__45234),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_14_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_14_27_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_14_27_6  (
            .in0(N__40801),
            .in1(N__45220),
            .in2(N__38929),
            .in3(N__44985),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_14_28_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_14_28_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_14_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42502),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49868),
            .ce(),
            .sr(N__49518));
    defparam CONSTANT_ONE_LUT4_LC_14_30_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_30_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_30_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_15_5_0  (
            .in0(N__43739),
            .in1(N__43723),
            .in2(_gnd_net_),
            .in3(N__48331),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50010),
            .ce(N__45824),
            .sr(N__49376));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_15_5_5  (
            .in0(N__48330),
            .in1(N__44087),
            .in2(_gnd_net_),
            .in3(N__44070),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50010),
            .ce(N__45824),
            .sr(N__49376));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_15_6_0  (
            .in0(N__43564),
            .in1(N__43187),
            .in2(_gnd_net_),
            .in3(N__48350),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__45827),
            .sr(N__49378));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_15_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_15_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_15_6_4  (
            .in0(N__47358),
            .in1(N__47387),
            .in2(_gnd_net_),
            .in3(N__48351),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__45827),
            .sr(N__49378));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_15_6_5  (
            .in0(N__48349),
            .in1(N__43205),
            .in2(_gnd_net_),
            .in3(N__43597),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__45827),
            .sr(N__49378));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_7_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_7_0  (
            .in0(N__39636),
            .in1(N__38901),
            .in2(N__39613),
            .in3(N__38938),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_15_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_15_7_1 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_15_7_1  (
            .in0(N__38937),
            .in1(N__39637),
            .in2(N__38905),
            .in3(N__39612),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_15_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_15_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_15_7_2  (
            .in0(N__47386),
            .in1(N__43660),
            .in2(N__47693),
            .in3(N__47323),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_15_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_15_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_15_7_4  (
            .in0(N__47594),
            .in1(N__41878),
            .in2(N__48623),
            .in3(N__41485),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_15_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_15_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_15_7_5  (
            .in0(N__45399),
            .in1(N__45369),
            .in2(_gnd_net_),
            .in3(N__48319),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_15_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_15_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_15_7_7  (
            .in0(N__43706),
            .in1(N__47224),
            .in2(N__47180),
            .in3(N__43846),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_15_8_0  (
            .in0(N__48324),
            .in1(N__43801),
            .in2(_gnd_net_),
            .in3(N__43771),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_1  (
            .in0(N__45537),
            .in1(N__45502),
            .in2(_gnd_net_),
            .in3(N__48326),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_15_8_2  (
            .in0(N__48323),
            .in1(N__45901),
            .in2(_gnd_net_),
            .in3(N__45928),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_15_8_3  (
            .in0(N__45397),
            .in1(N__45365),
            .in2(_gnd_net_),
            .in3(N__48327),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_15_8_4  (
            .in0(N__48322),
            .in1(N__45467),
            .in2(_gnd_net_),
            .in3(N__45442),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_15_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_15_8_6  (
            .in0(N__48321),
            .in1(N__43690),
            .in2(_gnd_net_),
            .in3(N__43661),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_7  (
            .in0(N__43825),
            .in1(N__43853),
            .in2(_gnd_net_),
            .in3(N__48325),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(N__45826),
            .sr(N__49387));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__39037),
            .in2(N__41104),
            .in3(N__39408),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__40987),
            .in2(N__39031),
            .in3(N__39382),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__39013),
            .in2(N__39022),
            .in3(N__39364),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__39007),
            .in2(N__39001),
            .in3(N__39346),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__38989),
            .in2(N__38983),
            .in3(N__39328),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_9_5  (
            .in0(N__39310),
            .in1(N__38971),
            .in2(N__38965),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__38956),
            .in2(N__38947),
            .in3(N__39292),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__39157),
            .in2(N__39145),
            .in3(N__39274),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__39136),
            .in2(N__39127),
            .in3(N__39547),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__41116),
            .in2(N__39118),
            .in3(N__39529),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__39097),
            .in2(N__39109),
            .in3(N__39511),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__39091),
            .in2(N__41095),
            .in3(N__39493),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_10_4  (
            .in0(N__39475),
            .in1(N__39073),
            .in2(N__39085),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__41359),
            .in2(N__39067),
            .in3(N__39457),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__39058),
            .in2(N__39049),
            .in3(N__39436),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__40813),
            .in2(N__40876),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__40909),
            .in2(N__40981),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__40996),
            .in2(N__41083),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__39256),
            .in2(N__39247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__39232),
            .in2(N__39223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__39211),
            .in2(N__39202),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__39190),
            .in2(N__39184),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_15_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_15_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__39175),
            .in2(N__39169),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39415),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__41341),
            .in2(N__39412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_12_1  (
            .in0(N__45773),
            .in1(N__39381),
            .in2(_gnd_net_),
            .in3(N__39367),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_12_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_12_2  (
            .in0(N__45832),
            .in1(N__39363),
            .in2(N__41317),
            .in3(N__39349),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_12_3  (
            .in0(N__45774),
            .in1(N__39345),
            .in2(_gnd_net_),
            .in3(N__39331),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_12_4  (
            .in0(N__45833),
            .in1(N__39327),
            .in2(_gnd_net_),
            .in3(N__39313),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_12_5  (
            .in0(N__45775),
            .in1(N__39309),
            .in2(_gnd_net_),
            .in3(N__39295),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_15_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_15_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_15_12_6  (
            .in0(N__45834),
            .in1(N__39291),
            .in2(_gnd_net_),
            .in3(N__39277),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_7  (
            .in0(N__45776),
            .in1(N__39273),
            .in2(_gnd_net_),
            .in3(N__39259),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49946),
            .ce(),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_13_0  (
            .in0(N__45780),
            .in1(N__39546),
            .in2(_gnd_net_),
            .in3(N__39532),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_15_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_15_13_1  (
            .in0(N__45769),
            .in1(N__39528),
            .in2(_gnd_net_),
            .in3(N__39514),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_15_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_15_13_2  (
            .in0(N__45777),
            .in1(N__39510),
            .in2(_gnd_net_),
            .in3(N__39496),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_15_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_15_13_3  (
            .in0(N__45770),
            .in1(N__39492),
            .in2(_gnd_net_),
            .in3(N__39478),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_15_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_15_13_4  (
            .in0(N__45778),
            .in1(N__39474),
            .in2(_gnd_net_),
            .in3(N__39460),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_15_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_15_13_5  (
            .in0(N__45771),
            .in1(N__39453),
            .in2(_gnd_net_),
            .in3(N__39439),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_15_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_15_13_6  (
            .in0(N__45779),
            .in1(N__39435),
            .in2(_gnd_net_),
            .in3(N__39421),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_15_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_15_13_7  (
            .in0(N__45772),
            .in1(N__40848),
            .in2(_gnd_net_),
            .in3(N__39418),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49934),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_14_0  (
            .in0(N__45757),
            .in1(N__40827),
            .in2(_gnd_net_),
            .in3(N__39652),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_14_1  (
            .in0(N__45781),
            .in1(N__40938),
            .in2(_gnd_net_),
            .in3(N__39649),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_14_2  (
            .in0(N__45758),
            .in1(N__40962),
            .in2(_gnd_net_),
            .in3(N__39646),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_15_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_15_14_3  (
            .in0(N__45782),
            .in1(N__41024),
            .in2(_gnd_net_),
            .in3(N__39643),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_15_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_15_14_4  (
            .in0(N__45759),
            .in1(N__41049),
            .in2(_gnd_net_),
            .in3(N__39640),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_15_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_15_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_15_14_5  (
            .in0(N__45783),
            .in1(N__39630),
            .in2(_gnd_net_),
            .in3(N__39616),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_15_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_15_14_6  (
            .in0(N__45760),
            .in1(N__39603),
            .in2(_gnd_net_),
            .in3(N__39589),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_15_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_15_14_7  (
            .in0(N__45784),
            .in1(N__39586),
            .in2(_gnd_net_),
            .in3(N__39571),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49926),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_15_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_15_15_0  (
            .in0(N__45753),
            .in1(N__39566),
            .in2(_gnd_net_),
            .in3(N__39550),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_15_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_15_15_1  (
            .in0(N__45814),
            .in1(N__39822),
            .in2(_gnd_net_),
            .in3(N__39808),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_15_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_15_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_15_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_15_15_2  (
            .in0(N__45754),
            .in1(N__39792),
            .in2(_gnd_net_),
            .in3(N__39778),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_15_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_15_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_15_15_3  (
            .in0(N__45815),
            .in1(N__39765),
            .in2(_gnd_net_),
            .in3(N__39751),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_15_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_15_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_15_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_15_15_4  (
            .in0(N__45755),
            .in1(N__39741),
            .in2(_gnd_net_),
            .in3(N__39727),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_15_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_15_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_15_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_15_15_5  (
            .in0(N__45816),
            .in1(N__39713),
            .in2(_gnd_net_),
            .in3(N__39697),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_15_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_15_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_15_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_15_15_6  (
            .in0(N__45756),
            .in1(N__39680),
            .in2(_gnd_net_),
            .in3(N__39694),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_tr.running_LC_15_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_15_15_7 .LUT_INIT=16'b1111010001110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_15_15_7  (
            .in0(N__41801),
            .in1(N__41760),
            .in2(N__41818),
            .in3(N__41842),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49435));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_15_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_15_16_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_15_16_2  (
            .in0(N__40014),
            .in1(N__41678),
            .in2(N__40036),
            .in3(N__41617),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__41718),
            .in2(_gnd_net_),
            .in3(N__42423),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_15_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_15_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__40031),
            .in2(_gnd_net_),
            .in3(N__40013),
            .lcout(\phase_controller_inst1.state_RNIE87FZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_15_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_15_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39982),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_15_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_15_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__46696),
            .in2(_gnd_net_),
            .in3(N__39932),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_15_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_15_18_0  (
            .in0(N__40047),
            .in1(N__40200),
            .in2(N__40231),
            .in3(N__40071),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_15_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__39864),
            .in2(_gnd_net_),
            .in3(N__39883),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_15_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_15_18_2  (
            .in0(N__40171),
            .in1(N__39874),
            .in2(N__39886),
            .in3(N__40186),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_15_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_15_18_4  (
            .in0(N__39882),
            .in1(N__39853),
            .in2(N__39844),
            .in3(N__40216),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_15_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_15_18_5  (
            .in0(N__39873),
            .in1(N__39865),
            .in2(N__39856),
            .in3(N__40117),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_15_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_15_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__39852),
            .in2(_gnd_net_),
            .in3(N__39840),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_15_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_15_19_0  (
            .in0(N__40227),
            .in1(N__40212),
            .in2(N__40201),
            .in3(N__40179),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_19_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_19_1  (
            .in0(N__40180),
            .in1(_gnd_net_),
            .in2(N__40135),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_15_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_15_19_2  (
            .in0(N__41967),
            .in1(N__40167),
            .in2(N__40156),
            .in3(N__41913),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_15_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_15_19_3  (
            .in0(N__40153),
            .in1(N__40087),
            .in2(N__40147),
            .in3(N__40144),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_15_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_15_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_15_19_4  (
            .in0(N__40098),
            .in1(N__40131),
            .in2(N__40111),
            .in3(N__40123),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_15_19_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__41931),
            .in2(_gnd_net_),
            .in3(N__41949),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_15_19_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_15_19_6  (
            .in0(N__40107),
            .in1(N__40056),
            .in2(N__40099),
            .in3(N__40080),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_15_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_15_19_7  (
            .in0(N__40081),
            .in1(N__40072),
            .in2(N__40060),
            .in3(N__40048),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_15_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_15_20_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_15_20_3  (
            .in0(N__42046),
            .in1(N__40384),
            .in2(N__42009),
            .in3(N__40365),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49892),
            .ce(),
            .sr(N__49475));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_21_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_21_7  (
            .in0(N__40382),
            .in1(N__42555),
            .in2(N__40366),
            .in3(N__42484),
            .lcout(\phase_controller_inst2.start_timer_tr_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_15_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_15_23_7 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_15_23_7  (
            .in0(N__40330),
            .in1(N__43307),
            .in2(N__42252),
            .in3(N__40306),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__44899),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__40288),
            .in2(_gnd_net_),
            .in3(N__40273),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__40270),
            .in2(_gnd_net_),
            .in3(N__40255),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(N__40252),
            .in2(_gnd_net_),
            .in3(N__40240),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__42856),
            .in2(_gnd_net_),
            .in3(N__40237),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__40465),
            .in2(N__42811),
            .in3(N__40234),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(N__42760),
            .in2(N__40497),
            .in3(N__40792),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__40469),
            .in2(N__42718),
            .in3(N__40399),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_27_0  (
            .in0(_gnd_net_),
            .in1(N__42670),
            .in2(_gnd_net_),
            .in3(N__40387),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_27_1  (
            .in0(_gnd_net_),
            .in1(N__42625),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_27_2  (
            .in0(_gnd_net_),
            .in1(N__42583),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_27_3  (
            .in0(_gnd_net_),
            .in1(N__43132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_27_4  (
            .in0(_gnd_net_),
            .in1(N__43084),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_27_5  (
            .in0(_gnd_net_),
            .in1(N__43036),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_27_6  (
            .in0(_gnd_net_),
            .in1(N__43003),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_27_7  (
            .in0(_gnd_net_),
            .in1(N__42976),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_28_0  (
            .in0(_gnd_net_),
            .in1(N__42949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_28_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_28_1  (
            .in0(_gnd_net_),
            .in1(N__42922),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_28_2  (
            .in0(_gnd_net_),
            .in1(N__43369),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_28_3  (
            .in0(_gnd_net_),
            .in1(N__43276),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_28_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40804),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_5_6  (
            .in0(N__48320),
            .in1(N__43743),
            .in2(_gnd_net_),
            .in3(N__43722),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_16_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_16_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_16_6_5  (
            .in0(N__43207),
            .in1(N__43605),
            .in2(_gnd_net_),
            .in3(N__48156),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_16_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_16_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_16_6_7  (
            .in0(N__45450),
            .in1(N__43414),
            .in2(N__45943),
            .in3(N__43472),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_7_0  (
            .in0(N__45513),
            .in1(N__45578),
            .in2(N__43895),
            .in3(N__48421),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_7_1  (
            .in0(N__40903),
            .in1(N__40897),
            .in2(N__40891),
            .in3(N__40888),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_7_2  (
            .in0(N__43507),
            .in1(N__48155),
            .in2(_gnd_net_),
            .in3(N__43481),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_7_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_7_3  (
            .in0(N__46181),
            .in1(N__41444),
            .in2(_gnd_net_),
            .in3(N__40882),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_7_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_7_4  (
            .in0(N__40833),
            .in1(N__45871),
            .in2(N__40861),
            .in3(N__45855),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_7_5 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_7_5  (
            .in0(N__45870),
            .in1(N__40860),
            .in2(N__45859),
            .in3(N__40834),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_7_6  (
            .in0(N__45471),
            .in1(N__45446),
            .in2(_gnd_net_),
            .in3(N__48153),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_7_7  (
            .in0(N__48154),
            .in1(N__43189),
            .in2(_gnd_net_),
            .in3(N__43572),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_16_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_16_8_1  (
            .in0(N__47296),
            .in1(N__47334),
            .in2(_gnd_net_),
            .in3(N__48173),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__45825),
            .sr(N__49381));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_8_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_16_8_2  (
            .in0(N__43913),
            .in1(_gnd_net_),
            .in2(N__43896),
            .in3(N__48175),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__45825),
            .sr(N__49381));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_16_8_3  (
            .in0(N__44188),
            .in1(N__44223),
            .in2(_gnd_net_),
            .in3(N__48171),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__45825),
            .sr(N__49381));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_16_8_6  (
            .in0(N__43488),
            .in1(N__43505),
            .in2(_gnd_net_),
            .in3(N__48174),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__45825),
            .sr(N__49381));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_16_8_7  (
            .in0(N__44167),
            .in1(N__44131),
            .in2(_gnd_net_),
            .in3(N__48172),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__45825),
            .sr(N__49381));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_9_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_9_0  (
            .in0(N__41031),
            .in1(N__41008),
            .in2(N__41059),
            .in3(N__41068),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_9_1  (
            .in0(N__41067),
            .in1(N__41058),
            .in2(N__41035),
            .in3(N__41007),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_16_9_7  (
            .in0(N__48328),
            .in1(N__43453),
            .in2(_gnd_net_),
            .in3(N__43422),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49981),
            .ce(N__45823),
            .sr(N__49388));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_10_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_10_0  (
            .in0(N__40969),
            .in1(N__40944),
            .in2(N__40924),
            .in3(N__41353),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_10_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_10_1  (
            .in0(N__41352),
            .in1(N__40968),
            .in2(N__40948),
            .in3(N__40920),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_16_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_16_10_5  (
            .in0(N__48267),
            .in1(N__47189),
            .in2(_gnd_net_),
            .in3(N__47154),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_10_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_16_10_6  (
            .in0(N__47190),
            .in1(_gnd_net_),
            .in2(N__41362),
            .in3(N__48269),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49971),
            .ce(N__45797),
            .sr(N__49395));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_16_10_7  (
            .in0(N__48268),
            .in1(N__45613),
            .in2(_gnd_net_),
            .in3(N__45582),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49971),
            .ce(N__45797),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_11_3  (
            .in0(N__48318),
            .in1(N__41445),
            .in2(_gnd_net_),
            .in3(N__41405),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_16_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_16_11_4  (
            .in0(N__41516),
            .in1(N__41493),
            .in2(_gnd_net_),
            .in3(N__48317),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_16_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_16_11_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__41802),
            .in2(_gnd_net_),
            .in3(N__41834),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_11_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_11_6  (
            .in0(N__41765),
            .in1(_gnd_net_),
            .in2(N__41344),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_16_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__41766),
            .in2(_gnd_net_),
            .in3(N__41328),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__41308),
            .in2(_gnd_net_),
            .in3(N__42146),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_12_2 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_12_2  (
            .in0(N__41587),
            .in1(N__41557),
            .in2(N__41542),
            .in3(N__41537),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(),
            .sr(N__49407));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_16_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_16_12_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_16_12_3  (
            .in0(N__46975),
            .in1(N__47014),
            .in2(N__46030),
            .in3(N__46865),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(),
            .sr(N__49407));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_13_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_13_0  (
            .in0(N__46549),
            .in1(N__46569),
            .in2(N__41383),
            .in3(N__41455),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_13_1  (
            .in0(N__41454),
            .in1(N__46548),
            .in2(N__46573),
            .in3(N__41379),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_16_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_16_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_16_13_2  (
            .in0(N__41517),
            .in1(N__41494),
            .in2(_gnd_net_),
            .in3(N__48389),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__47916),
            .sr(N__49414));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_16_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_16_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_16_13_3  (
            .in0(N__48385),
            .in1(N__41446),
            .in2(_gnd_net_),
            .in3(N__41406),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__47916),
            .sr(N__49414));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_16_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_16_13_4  (
            .in0(N__46147),
            .in1(N__48390),
            .in2(_gnd_net_),
            .in3(N__46185),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__47916),
            .sr(N__49414));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_16_13_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_16_13_5  (
            .in0(N__41370),
            .in1(N__46498),
            .in2(N__46528),
            .in3(N__41850),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_16_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_16_13_6 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_16_13_6  (
            .in0(N__46524),
            .in1(N__46497),
            .in2(N__41854),
            .in3(N__41371),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_16_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_16_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_16_13_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__41902),
            .in2(N__48400),
            .in3(N__41884),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__47916),
            .sr(N__49414));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_16_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42093),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49935),
            .ce(),
            .sr(N__49420));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_14_6 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_16_14_6  (
            .in0(N__41646),
            .in1(N__41761),
            .in2(N__41803),
            .in3(N__41841),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49935),
            .ce(),
            .sr(N__49420));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_16_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_16_15_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__41794),
            .in2(_gnd_net_),
            .in3(N__42086),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_15_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_15_4  (
            .in0(N__41814),
            .in1(N__41793),
            .in2(_gnd_net_),
            .in3(N__42085),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__41642),
            .in2(_gnd_net_),
            .in3(N__41598),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_16_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_16_16_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.state_1_LC_16_16_1  (
            .in0(N__41619),
            .in1(N__41734),
            .in2(_gnd_net_),
            .in3(N__41680),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.state_3_LC_16_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_16_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_16_16_2 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst1.state_3_LC_16_16_2  (
            .in0(N__42435),
            .in1(N__41719),
            .in2(N__42118),
            .in3(N__44683),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.state_0_LC_16_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_16_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_16_16_4 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_0_LC_16_16_4  (
            .in0(N__41679),
            .in1(N__41599),
            .in2(N__41650),
            .in3(N__41618),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst2.start_timer_hc_LC_16_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_16_16_6 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_16_16_6  (
            .in0(N__44733),
            .in1(N__42523),
            .in2(N__42067),
            .in3(N__42140),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.start_timer_tr_LC_16_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_16_7 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_16_16_7  (
            .in0(N__42111),
            .in1(N__42100),
            .in2(N__42094),
            .in3(N__44734),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__42033),
            .in2(_gnd_net_),
            .in3(N__41989),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_16_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_16_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_16_18_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_0_LC_16_18_0  (
            .in0(N__42554),
            .in1(N__44671),
            .in2(N__42501),
            .in3(N__44659),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(),
            .sr(N__49454));
    defparam \phase_controller_inst1.state_4_LC_16_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_16_18_1 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_16_18_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__44795),
            .in2(_gnd_net_),
            .in3(N__44729),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(),
            .sr(N__49454));
    defparam \phase_controller_inst2.start_timer_tr_LC_16_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_16_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_16_18_4 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_16_18_4  (
            .in0(N__44728),
            .in1(N__42058),
            .in2(N__46939),
            .in3(N__44638),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(),
            .sr(N__49454));
    defparam \phase_controller_inst2.state_3_LC_16_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_16_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_16_18_6 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_16_18_6  (
            .in0(N__42045),
            .in1(N__44682),
            .in2(N__42005),
            .in3(N__44637),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(),
            .sr(N__49454));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_19_2  (
            .in0(N__41971),
            .in1(N__41953),
            .in2(N__41938),
            .in3(N__41920),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_19_3  (
            .in0(N__42577),
            .in1(N__42571),
            .in2(N__42565),
            .in3(N__42562),
            .lcout(\current_shift_inst.PI_CTRL.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_16_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_16_21_4 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_16_21_4  (
            .in0(N__42556),
            .in1(N__42491),
            .in2(_gnd_net_),
            .in3(N__42516),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49893),
            .ce(),
            .sr(N__49476));
    defparam \phase_controller_inst1.test22_LC_16_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.test22_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test22_LC_16_21_7 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \phase_controller_inst1.test22_LC_16_21_7  (
            .in0(N__42387),
            .in1(N__42436),
            .in2(N__44740),
            .in3(N__44804),
            .lcout(test22_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49893),
            .ce(),
            .sr(N__49476));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_16_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50241),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(),
            .sr(N__49486));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_26_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_26_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_26_0  (
            .in0(_gnd_net_),
            .in1(N__42192),
            .in2(_gnd_net_),
            .in3(N__44844),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_16_26_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_16_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_16_26_1  (
            .in0(N__45268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42180),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2  (
            .in0(N__42181),
            .in1(N__45256),
            .in2(N__42172),
            .in3(N__44971),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5  (
            .in0(_gnd_net_),
            .in1(N__45300),
            .in2(_gnd_net_),
            .in3(N__42159),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_26_6  (
            .in0(N__45200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43242),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_7  (
            .in0(_gnd_net_),
            .in1(N__42909),
            .in2(_gnd_net_),
            .in3(N__45336),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_27_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_16_27_0  (
            .in0(_gnd_net_),
            .in1(N__42898),
            .in2(N__42877),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_16_27_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_27_1  (
            .in0(_gnd_net_),
            .in1(N__42850),
            .in2(N__42832),
            .in3(N__42802),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_27_2  (
            .in0(_gnd_net_),
            .in1(N__42799),
            .in2(N__42781),
            .in3(N__42754),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(N__42751),
            .in2(N__42733),
            .in3(N__42709),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_27_4  (
            .in0(_gnd_net_),
            .in1(N__42706),
            .in2(N__42691),
            .in3(N__42664),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_27_5  (
            .in0(_gnd_net_),
            .in1(N__42661),
            .in2(N__42643),
            .in3(N__42619),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_27_6  (
            .in0(_gnd_net_),
            .in1(N__42616),
            .in2(N__42604),
            .in3(N__43171),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_27_7  (
            .in0(_gnd_net_),
            .in1(N__43168),
            .in2(N__43153),
            .in3(N__43126),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_28_0  (
            .in0(_gnd_net_),
            .in1(N__43123),
            .in2(N__43108),
            .in3(N__43078),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_16_28_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_28_1  (
            .in0(_gnd_net_),
            .in1(N__43075),
            .in2(N__43057),
            .in3(N__43030),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_28_2  (
            .in0(_gnd_net_),
            .in1(N__43327),
            .in2(N__43027),
            .in3(N__42997),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_28_3  (
            .in0(_gnd_net_),
            .in1(N__42994),
            .in2(N__43340),
            .in3(N__42970),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_28_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_28_4  (
            .in0(_gnd_net_),
            .in1(N__43331),
            .in2(N__42967),
            .in3(N__42943),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_28_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_28_5  (
            .in0(_gnd_net_),
            .in1(N__42940),
            .in2(N__43341),
            .in3(N__42916),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_28_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_28_6  (
            .in0(_gnd_net_),
            .in1(N__43335),
            .in2(N__43390),
            .in3(N__43363),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_28_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_28_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_28_7  (
            .in0(_gnd_net_),
            .in1(N__43360),
            .in2(N__43342),
            .in3(N__43270),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_29_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_29_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_29_0  (
            .in0(N__43267),
            .in1(N__43261),
            .in2(_gnd_net_),
            .in3(N__43249),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_16_29_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_16_29_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_16_29_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_16_29_2  (
            .in0(N__43246),
            .in1(N__45201),
            .in2(N__44972),
            .in3(N__45178),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_16_29_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_16_29_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_16_29_4 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_16_29_4  (
            .in0(N__44945),
            .in1(N__45130),
            .in2(N__45154),
            .in3(N__45247),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_17_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_17_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_17_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_17_6_3  (
            .in0(N__43206),
            .in1(N__43606),
            .in2(_gnd_net_),
            .in3(N__48170),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__47911),
            .sr(N__49374));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_17_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_17_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_17_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_17_6_5  (
            .in0(N__43188),
            .in1(N__43573),
            .in2(_gnd_net_),
            .in3(N__48169),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__47911),
            .sr(N__49374));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_17_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_17_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_17_7_0  (
            .in0(N__43821),
            .in1(N__43858),
            .in2(_gnd_net_),
            .in3(N__48221),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_7_1  (
            .in0(N__48223),
            .in1(N__43915),
            .in2(_gnd_net_),
            .in3(N__43888),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(N__43990),
            .in2(_gnd_net_),
            .in3(N__44065),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_7_3  (
            .in0(N__48222),
            .in1(N__43689),
            .in2(_gnd_net_),
            .in3(N__43662),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_17_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_17_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_17_7_4  (
            .in0(N__43598),
            .in1(N__43565),
            .in2(N__44137),
            .in3(N__44215),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5  (
            .in0(N__45398),
            .in1(N__43772),
            .in2(N__43534),
            .in3(N__43531),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_6  (
            .in0(N__47543),
            .in1(N__43525),
            .in2(N__43519),
            .in3(N__43516),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_17_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_17_7_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_17_7_7  (
            .in0(N__44216),
            .in1(_gnd_net_),
            .in2(N__43510),
            .in3(N__44186),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_17_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_17_8_0  (
            .in0(N__48157),
            .in1(N__43506),
            .in2(_gnd_net_),
            .in3(N__43489),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_17_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_17_8_1  (
            .in0(N__45900),
            .in1(N__45941),
            .in2(_gnd_net_),
            .in3(N__48163),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_17_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_17_8_2  (
            .in0(N__48159),
            .in1(N__43449),
            .in2(_gnd_net_),
            .in3(N__43426),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_17_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_17_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_17_8_3  (
            .in0(N__47292),
            .in1(N__47335),
            .in2(_gnd_net_),
            .in3(N__48162),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_17_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_17_8_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_17_8_4  (
            .in0(N__48158),
            .in1(N__43914),
            .in2(N__43897),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_17_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_17_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_17_8_5  (
            .in0(N__43857),
            .in1(N__43817),
            .in2(_gnd_net_),
            .in3(N__48160),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_6  (
            .in0(N__43800),
            .in1(N__48164),
            .in2(_gnd_net_),
            .in3(N__43780),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_17_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_17_8_7  (
            .in0(N__43744),
            .in1(N__43721),
            .in2(_gnd_net_),
            .in3(N__48161),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__47912),
            .sr(N__49379));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_9_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_9_0  (
            .in0(N__46626),
            .in1(N__46605),
            .in2(N__43618),
            .in3(N__43627),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_17_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_17_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_17_9_1  (
            .in0(N__43626),
            .in1(N__46627),
            .in2(N__46606),
            .in3(N__43614),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_17_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_17_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_17_9_2  (
            .in0(N__48270),
            .in1(N__43685),
            .in2(_gnd_net_),
            .in3(N__43663),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49994),
            .ce(N__47913),
            .sr(N__49382));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_17_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_17_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_17_9_3  (
            .in0(N__47362),
            .in1(N__47397),
            .in2(_gnd_net_),
            .in3(N__48273),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49994),
            .ce(N__47913),
            .sr(N__49382));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_17_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_17_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_17_9_5  (
            .in0(N__44224),
            .in1(N__44187),
            .in2(_gnd_net_),
            .in3(N__48271),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49994),
            .ce(N__47913),
            .sr(N__49382));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_17_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_17_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_17_9_7  (
            .in0(N__44163),
            .in1(N__44136),
            .in2(_gnd_net_),
            .in3(N__48272),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49994),
            .ce(N__47913),
            .sr(N__49382));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0  (
            .in0(N__46098),
            .in1(N__46336),
            .in2(N__46363),
            .in3(N__46114),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_17_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_17_10_5  (
            .in0(N__44098),
            .in1(N__44071),
            .in2(_gnd_net_),
            .in3(N__48275),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49982),
            .ce(N__47915),
            .sr(N__49389));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_17_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_17_10_6  (
            .in0(N__44034),
            .in1(N__48274),
            .in2(_gnd_net_),
            .in3(N__44002),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49982),
            .ce(N__47915),
            .sr(N__49389));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_17_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_17_11_0  (
            .in0(N__46016),
            .in1(N__43945),
            .in2(N__43960),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_17_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__43927),
            .in2(N__43939),
            .in3(N__46002),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_17_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__43921),
            .in2(N__45415),
            .in3(N__45972),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_17_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_17_11_3  (
            .in0(N__45957),
            .in1(N__44371),
            .in2(N__44359),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_17_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__45349),
            .in2(N__44347),
            .in3(N__46311),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_17_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_17_11_5  (
            .in0(N__46297),
            .in1(N__44338),
            .in2(N__44329),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_17_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__44320),
            .in2(N__44314),
            .in3(N__46278),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_17_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__44305),
            .in2(N__44299),
            .in3(N__46264),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_17_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__44287),
            .in2(N__44278),
            .in3(N__46245),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_17_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__44269),
            .in2(N__44260),
            .in3(N__46230),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_17_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_17_12_2  (
            .in0(N__46215),
            .in1(N__44248),
            .in2(N__44236),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_17_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_17_12_3  (
            .in0(N__46200),
            .in1(N__44452),
            .in2(N__44464),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_17_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__44434),
            .in2(N__44446),
            .in3(N__46473),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_17_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_17_12_5  (
            .in0(N__46458),
            .in1(N__47143),
            .in2(N__44428),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_17_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_17_12_6  (
            .in0(N__46443),
            .in1(N__44419),
            .in2(N__44410),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_17_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_17_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__47206),
            .in2(N__47059),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_17_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_17_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__46042),
            .in2(N__45628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_17_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_17_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__44401),
            .in2(N__46081),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_17_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_17_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__44392),
            .in2(N__44383),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_17_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_17_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__47734),
            .in2(N__47794),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_17_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_17_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__44524),
            .in2(N__44518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_17_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_17_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__44509),
            .in2(N__44503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_17_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_17_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__47470),
            .in2(N__47410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_17_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_17_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44494),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_17_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_17_14_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__46902),
            .in2(_gnd_net_),
            .in3(N__47030),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_17_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_17_14_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44491),
            .in3(N__46967),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_17_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_17_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_17_15_3  (
            .in0(N__46942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(),
            .sr(N__49421));
    defparam \phase_controller_inst1.test_LC_17_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.test_LC_17_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test_LC_17_16_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \phase_controller_inst1.test_LC_17_16_3  (
            .in0(N__44475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44735),
            .lcout(test_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(),
            .sr(N__49429));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_16_7 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_17_16_7  (
            .in0(N__44657),
            .in1(N__46968),
            .in2(N__46911),
            .in3(N__47035),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(),
            .sr(N__49429));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__44777),
            .in2(_gnd_net_),
            .in3(N__44713),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_17_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_17_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__44670),
            .in2(_gnd_net_),
            .in3(N__44658),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_17_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_17_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__44611),
            .in2(_gnd_net_),
            .in3(N__44629),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_17_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_17_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__44587),
            .in2(_gnd_net_),
            .in3(N__44605),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_17_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_17_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_17_26_2  (
            .in0(_gnd_net_),
            .in1(N__44566),
            .in2(_gnd_net_),
            .in3(N__44581),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_17_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_17_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_17_26_3  (
            .in0(_gnd_net_),
            .in1(N__44548),
            .in2(_gnd_net_),
            .in3(N__44560),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_17_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_17_26_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__44530),
            .in2(_gnd_net_),
            .in3(N__44542),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_17_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_17_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_17_26_5  (
            .in0(_gnd_net_),
            .in1(N__45100),
            .in2(_gnd_net_),
            .in3(N__45115),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_17_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_17_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_17_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_17_26_6  (
            .in0(_gnd_net_),
            .in1(N__45079),
            .in2(_gnd_net_),
            .in3(N__45094),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_17_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_17_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_17_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_17_26_7  (
            .in0(_gnd_net_),
            .in1(N__45058),
            .in2(_gnd_net_),
            .in3(N__45073),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_17_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_17_27_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__45034),
            .in2(_gnd_net_),
            .in3(N__45052),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_17_27_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_17_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_17_27_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_17_27_1  (
            .in0(_gnd_net_),
            .in1(N__45010),
            .in2(_gnd_net_),
            .in3(N__45028),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_17_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_17_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_17_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_17_27_2  (
            .in0(_gnd_net_),
            .in1(N__46649),
            .in2(_gnd_net_),
            .in3(N__44995),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_17_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_17_27_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_17_27_3  (
            .in0(N__44949),
            .in1(N__44898),
            .in2(_gnd_net_),
            .in3(N__44854),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_17_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_17_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_17_27_4  (
            .in0(_gnd_net_),
            .in1(N__44840),
            .in2(_gnd_net_),
            .in3(N__44815),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_17_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_17_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_17_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_17_27_5  (
            .in0(_gnd_net_),
            .in1(N__45332),
            .in2(_gnd_net_),
            .in3(N__45307),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_17_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_17_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_17_27_6  (
            .in0(_gnd_net_),
            .in1(N__45296),
            .in2(_gnd_net_),
            .in3(N__45271),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_17_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_17_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_17_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_17_27_7  (
            .in0(_gnd_net_),
            .in1(N__45267),
            .in2(_gnd_net_),
            .in3(N__45250),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_17_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_17_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_17_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_17_28_0  (
            .in0(_gnd_net_),
            .in1(N__45128),
            .in2(_gnd_net_),
            .in3(N__45241),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_17_28_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_17_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_17_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_17_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_17_28_1  (
            .in0(_gnd_net_),
            .in1(N__45238),
            .in2(_gnd_net_),
            .in3(N__45205),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_17_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_17_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_17_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_17_28_2  (
            .in0(_gnd_net_),
            .in1(N__45202),
            .in2(_gnd_net_),
            .in3(N__45172),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_17_28_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_17_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_17_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_17_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45169),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_17_28_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_17_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_17_28_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_17_28_5  (
            .in0(N__45129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45153),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_5_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_5_0  (
            .in0(N__45893),
            .in1(N__45942),
            .in2(_gnd_net_),
            .in3(N__48276),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_6_2  (
            .in0(N__45605),
            .in1(N__45583),
            .in2(_gnd_net_),
            .in3(N__48152),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_18_7_1  (
            .in0(N__47271),
            .in1(N__47244),
            .in2(_gnd_net_),
            .in3(N__48242),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50016),
            .ce(N__45836),
            .sr(N__49375));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_18_7_7  (
            .in0(N__48459),
            .in1(N__48432),
            .in2(_gnd_net_),
            .in3(N__48243),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50016),
            .ce(N__45836),
            .sr(N__49375));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_18_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_18_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_18_8_1  (
            .in0(N__46065),
            .in1(N__46419),
            .in2(N__46393),
            .in3(N__46053),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_18_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_18_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_18_8_2  (
            .in0(N__45606),
            .in1(N__45574),
            .in2(_gnd_net_),
            .in3(N__48168),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(N__47914),
            .sr(N__49377));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_18_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_18_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_18_8_3  (
            .in0(N__48165),
            .in1(N__45541),
            .in2(_gnd_net_),
            .in3(N__45514),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(N__47914),
            .sr(N__49377));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_18_8_5  (
            .in0(N__48166),
            .in1(N__45475),
            .in2(_gnd_net_),
            .in3(N__45451),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(N__47914),
            .sr(N__49377));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_18_8_7  (
            .in0(N__48167),
            .in1(N__45403),
            .in2(_gnd_net_),
            .in3(N__45373),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(N__47914),
            .sr(N__49377));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_9_1  (
            .in0(N__48277),
            .in1(N__46186),
            .in2(_gnd_net_),
            .in3(N__46136),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_5 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_5  (
            .in0(N__46110),
            .in1(N__46335),
            .in2(N__46099),
            .in3(N__46359),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_9_6  (
            .in0(N__47270),
            .in1(N__47243),
            .in2(_gnd_net_),
            .in3(N__48278),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_9_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_9_7  (
            .in0(N__46066),
            .in1(N__46392),
            .in2(N__46423),
            .in3(N__46054),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__46029),
            .in2(N__46999),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_10_1  (
            .in0(N__46824),
            .in1(N__46003),
            .in2(_gnd_net_),
            .in3(N__45991),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_10_2  (
            .in0(N__46866),
            .in1(N__45988),
            .in2(N__45976),
            .in3(N__45961),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_10_3  (
            .in0(N__46825),
            .in1(N__45958),
            .in2(_gnd_net_),
            .in3(N__45946),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_10_4  (
            .in0(N__46867),
            .in1(N__46312),
            .in2(_gnd_net_),
            .in3(N__46300),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_10_5  (
            .in0(N__46826),
            .in1(N__46296),
            .in2(_gnd_net_),
            .in3(N__46282),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_10_6  (
            .in0(N__46868),
            .in1(N__46279),
            .in2(_gnd_net_),
            .in3(N__46267),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_10_7  (
            .in0(N__46827),
            .in1(N__46263),
            .in2(_gnd_net_),
            .in3(N__46249),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49995),
            .ce(),
            .sr(N__49383));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_11_0  (
            .in0(N__46835),
            .in1(N__46246),
            .in2(_gnd_net_),
            .in3(N__46234),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_11_1  (
            .in0(N__46820),
            .in1(N__46231),
            .in2(_gnd_net_),
            .in3(N__46219),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_11_2  (
            .in0(N__46832),
            .in1(N__46216),
            .in2(_gnd_net_),
            .in3(N__46204),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_11_3  (
            .in0(N__46821),
            .in1(N__46201),
            .in2(_gnd_net_),
            .in3(N__46189),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_11_4  (
            .in0(N__46833),
            .in1(N__46474),
            .in2(_gnd_net_),
            .in3(N__46462),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_11_5  (
            .in0(N__46822),
            .in1(N__46459),
            .in2(_gnd_net_),
            .in3(N__46447),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_11_6  (
            .in0(N__46834),
            .in1(N__46444),
            .in2(_gnd_net_),
            .in3(N__46432),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_11_7  (
            .in0(N__46823),
            .in1(N__47078),
            .in2(_gnd_net_),
            .in3(N__46429),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49983),
            .ce(),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_12_0  (
            .in0(N__46828),
            .in1(N__47126),
            .in2(_gnd_net_),
            .in3(N__46426),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_12_1  (
            .in0(N__46869),
            .in1(N__46418),
            .in2(_gnd_net_),
            .in3(N__46396),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_12_2  (
            .in0(N__46829),
            .in1(N__46388),
            .in2(_gnd_net_),
            .in3(N__46366),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_18_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_18_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_18_12_3  (
            .in0(N__46870),
            .in1(N__46358),
            .in2(_gnd_net_),
            .in3(N__46339),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_18_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_18_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_18_12_4  (
            .in0(N__46830),
            .in1(N__46334),
            .in2(_gnd_net_),
            .in3(N__46315),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_18_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_18_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_18_12_5  (
            .in0(N__46871),
            .in1(N__46625),
            .in2(_gnd_net_),
            .in3(N__46609),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_18_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_18_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_18_12_6  (
            .in0(N__46831),
            .in1(N__46596),
            .in2(_gnd_net_),
            .in3(N__46582),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_18_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_18_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_18_12_7  (
            .in0(N__46872),
            .in1(N__47769),
            .in2(_gnd_net_),
            .in3(N__46579),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49972),
            .ce(),
            .sr(N__49396));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_18_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_18_13_0  (
            .in0(N__46842),
            .in1(N__47754),
            .in2(_gnd_net_),
            .in3(N__46576),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_18_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_18_13_1  (
            .in0(N__46836),
            .in1(N__46568),
            .in2(_gnd_net_),
            .in3(N__46552),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_18_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_18_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_18_13_2  (
            .in0(N__46843),
            .in1(N__46547),
            .in2(_gnd_net_),
            .in3(N__46531),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_18_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_18_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_18_13_3  (
            .in0(N__46837),
            .in1(N__46523),
            .in2(_gnd_net_),
            .in3(N__46501),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_18_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_18_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_18_13_4  (
            .in0(N__46844),
            .in1(N__46496),
            .in2(_gnd_net_),
            .in3(N__46477),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_18_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_18_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_18_13_5  (
            .in0(N__46838),
            .in1(N__47447),
            .in2(_gnd_net_),
            .in3(N__47041),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_18_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_18_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_18_13_6  (
            .in0(N__46845),
            .in1(N__47426),
            .in2(_gnd_net_),
            .in3(N__47038),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49962),
            .ce(),
            .sr(N__49401));
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_14_3 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_18_14_3  (
            .in0(N__46987),
            .in1(N__46966),
            .in2(N__46912),
            .in3(N__47034),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(),
            .sr(N__49408));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__46965),
            .in2(_gnd_net_),
            .in3(N__47010),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_15_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_15_2  (
            .in0(N__46903),
            .in1(N__46986),
            .in2(_gnd_net_),
            .in3(N__46940),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_18_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_18_15_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_18_15_3  (
            .in0(N__46941),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46904),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46726),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49422));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_18_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_18_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_18_27_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_18_27_6  (
            .in0(_gnd_net_),
            .in1(N__46674),
            .in2(_gnd_net_),
            .in3(N__46653),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50023),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_6_5  (
            .in0(N__47357),
            .in1(N__47398),
            .in2(_gnd_net_),
            .in3(N__48315),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_20_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_20_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_20_8_5  (
            .in0(N__47291),
            .in1(N__47333),
            .in2(_gnd_net_),
            .in3(N__48297),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_20_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_20_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_20_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_20_9_7  (
            .in0(N__48298),
            .in1(N__47272),
            .in2(_gnd_net_),
            .in3(N__47248),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50017),
            .ce(N__47917),
            .sr(N__49380));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_20_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_20_10_0 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_20_10_0  (
            .in0(N__47932),
            .in1(N__47103),
            .in2(N__47131),
            .in3(N__47088),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_20_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_20_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_20_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_20_10_5  (
            .in0(N__48299),
            .in1(N__47194),
            .in2(_gnd_net_),
            .in3(N__47158),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50012),
            .ce(N__47918),
            .sr(N__49384));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_20_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_20_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_20_11_1  (
            .in0(N__47492),
            .in1(N__47544),
            .in2(_gnd_net_),
            .in3(N__48282),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_20_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_20_11_3 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_20_11_3  (
            .in0(N__47127),
            .in1(N__47104),
            .in2(N__47089),
            .in3(N__47931),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_4  (
            .in0(N__48283),
            .in1(N__47624),
            .in2(_gnd_net_),
            .in3(N__47601),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_20_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_20_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_20_11_7  (
            .in0(N__48647),
            .in1(N__48624),
            .in2(_gnd_net_),
            .in3(N__48284),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_20_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_20_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_20_12_3  (
            .in0(N__47715),
            .in1(N__47694),
            .in2(_gnd_net_),
            .in3(N__48353),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_13_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_13_0  (
            .in0(N__47554),
            .in1(N__47641),
            .in2(N__47779),
            .in3(N__47753),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_13_1  (
            .in0(N__47640),
            .in1(N__47775),
            .in2(N__47755),
            .in3(N__47553),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_20_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_20_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_20_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_20_13_2  (
            .in0(N__48354),
            .in1(N__47711),
            .in2(_gnd_net_),
            .in3(N__47695),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__47920),
            .sr(N__49402));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_20_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_20_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_20_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_20_13_3  (
            .in0(N__47625),
            .in1(N__47602),
            .in2(_gnd_net_),
            .in3(N__48356),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__47920),
            .sr(N__49402));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_20_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_20_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_20_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_20_13_4  (
            .in0(N__48355),
            .in1(N__47545),
            .in2(_gnd_net_),
            .in3(N__47496),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__47920),
            .sr(N__49402));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_20_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_20_13_5 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_20_13_5  (
            .in0(N__48579),
            .in1(N__47451),
            .in2(N__47431),
            .in3(N__47460),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_20_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_20_13_6 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_20_13_6  (
            .in0(N__47461),
            .in1(N__48580),
            .in2(N__47452),
            .in3(N__47430),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_20_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_20_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_20_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_20_13_7  (
            .in0(N__48648),
            .in1(N__48625),
            .in2(_gnd_net_),
            .in3(N__48357),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__47920),
            .sr(N__49402));
    defparam \delay_measurement_inst.stop_timer_tr_LC_20_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_20_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_20_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48494),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(),
            .sr(N__49437));
    defparam \delay_measurement_inst.start_timer_tr_LC_20_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_20_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_20_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48493),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(),
            .sr(N__49437));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_21_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_21_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_21_7_0  (
            .in0(N__48458),
            .in1(N__48431),
            .in2(_gnd_net_),
            .in3(N__48316),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_21_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_21_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_21_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_21_10_4  (
            .in0(N__48460),
            .in1(N__48436),
            .in2(_gnd_net_),
            .in3(N__48352),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50018),
            .ce(N__47919),
            .sr(N__49391));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_21_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_21_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_21_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47884),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_22_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_22_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_22_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_22_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47860),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49482));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_7 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_7  (
            .in0(N__48667),
            .in1(N__48721),
            .in2(N__48880),
            .in3(N__48661),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_20_1  (
            .in0(_gnd_net_),
            .in1(N__48897),
            .in2(_gnd_net_),
            .in3(N__48773),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_20_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_20_2  (
            .in0(_gnd_net_),
            .in1(N__50405),
            .in2(_gnd_net_),
            .in3(N__50297),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_20_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_20_3  (
            .in0(N__50345),
            .in1(N__50505),
            .in2(N__48691),
            .in3(N__50178),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_21_2 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_21_2  (
            .in0(N__50243),
            .in1(N__48683),
            .in2(N__48923),
            .in3(N__50123),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_21_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_21_6  (
            .in0(N__50242),
            .in1(N__48684),
            .in2(_gnd_net_),
            .in3(N__50122),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_5  (
            .in0(N__50244),
            .in1(N__48688),
            .in2(N__48924),
            .in3(N__50124),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_1  (
            .in0(_gnd_net_),
            .in1(N__50468),
            .in2(_gnd_net_),
            .in3(N__50264),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_2  (
            .in0(N__50321),
            .in1(N__50375),
            .in2(N__48670),
            .in3(N__50039),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_5  (
            .in0(N__50430),
            .in1(N__48954),
            .in2(_gnd_net_),
            .in3(N__48819),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_6  (
            .in0(N__50322),
            .in1(N__50376),
            .in2(N__50473),
            .in3(N__50040),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_24_2 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_24_2  (
            .in0(N__48655),
            .in1(N__48720),
            .in2(N__48876),
            .in3(N__50265),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_24_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_24_20_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_24_20_0  (
            .in0(N__50174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50412),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_24_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_24_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_24_20_1  (
            .in0(N__50298),
            .in1(N__50352),
            .in2(N__48997),
            .in3(N__50501),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_20_2 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_20_2  (
            .in0(N__50240),
            .in1(N__48994),
            .in2(N__48988),
            .in3(N__50063),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_21_0 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_21_0  (
            .in0(N__48786),
            .in1(N__48798),
            .in2(N__48985),
            .in3(N__48774),
            .lcout(\current_shift_inst.PI_CTRL.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_0  (
            .in0(_gnd_net_),
            .in1(N__48976),
            .in2(_gnd_net_),
            .in3(N__50443),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_1 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_1  (
            .in0(N__48940),
            .in1(N__48931),
            .in2(N__48925),
            .in3(N__50079),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_2  (
            .in0(_gnd_net_),
            .in1(N__48841),
            .in2(_gnd_net_),
            .in3(N__50442),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_4  (
            .in0(N__48805),
            .in1(N__48787),
            .in2(_gnd_net_),
            .in3(N__48775),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_5 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_5  (
            .in0(N__50245),
            .in1(N__50121),
            .in2(N__50506),
            .in3(N__50078),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_6  (
            .in0(N__50452),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50441),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49490));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_1 .LUT_INIT=16'b1101110001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_1  (
            .in0(N__50239),
            .in1(N__50416),
            .in2(N__50143),
            .in3(N__50083),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49494));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_2 .LUT_INIT=16'b1011001110110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_2  (
            .in0(N__50082),
            .in1(N__50238),
            .in2(N__50359),
            .in3(N__50141),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49494));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_6 .LUT_INIT=16'b1011001110110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_6  (
            .in0(N__50080),
            .in1(N__50236),
            .in2(N__50305),
            .in3(N__50140),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49494));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_7 .LUT_INIT=16'b1101110001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_7  (
            .in0(N__50237),
            .in1(N__50179),
            .in2(N__50142),
            .in3(N__50081),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49494));
endmodule // MAIN
