-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Nov 29 2024 16:50:30

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    test : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    test22 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50662\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal un7_start_stop_0_a3 : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \N_39_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.timer_s1.N_161_i\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_199_i\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_198_i\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_8_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.N_1306_i\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal s1_phy_c : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal s3_phy_c : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.N_161_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \bfn_12_26_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \GB_BUFFER_red_c_g_THRU_CO\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_201_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal s2_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \bfn_13_27_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_200_i\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.state_RNIE87FZ0Z_2\ : std_logic;
signal il_max_comp1_c : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal state_3 : std_logic;
signal test22_c : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_16_27_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_16_28_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_16_29_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal test_c : std_logic;
signal start_stop_c : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_17_27_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_17_28_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_160\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_158\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clock_output_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal test_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal test22_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    test <= test_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    test22 <= test22_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__21079\&\N__34210\&\N__35644\&\N__21052\&\N__21007\&\N__21193\&\N__34330\&\N__29926\&\N__34177\&\N__34021\&\N__34243\&\N__33960\&\N__34354\&\N__34273\&\N__33937\&\N__21034\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40579\&'0'&\N__40578\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__42374\&\N__42367\&\N__42372\&\N__42366\&\N__42373\&\N__42365\&\N__42375\&\N__42362\&\N__42368\&\N__42361\&\N__42369\&\N__42363\&\N__42370\&\N__42364\&\N__42371\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40611\&\N__40608\&'0'&'0'&'0'&\N__40606\&\N__40610\&\N__40607\&\N__40609\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__42351\&\N__42354\&\N__42352\&\N__42355\&\N__42353\&\N__50377\&\N__50323\&\N__50472\&\N__50041\&\N__50266\&\N__48875\&\N__48716\&\N__48958\&\N__48823\&\N__50431\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40575\&\N__40572\&'0'&'0'&'0'&\N__40570\&\N__40574\&\N__40571\&\N__40573\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__34383\&\N__34299\&\N__36684\&\N__29980\&\N__36742\&\N__34407\&\N__34047\&\N__31029\&\N__36714\&\N__39981\&\N__34077\&\N__33993\&\N__29949\&\N__46722\&\N__47880\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__40787\&'0'&\N__40786\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__28675\,
            RESETB => \N__33031\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40789\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40577\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40655\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40605\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40576\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40569\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__40788\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__40782\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50660\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50662\,
            DIN => \N__50661\,
            DOUT => \N__50660\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50662\,
            PADOUT => \N__50661\,
            PADIN => \N__50660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50651\,
            DIN => \N__50650\,
            DOUT => \N__50649\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50651\,
            PADOUT => \N__50650\,
            PADIN => \N__50649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__46633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50642\,
            DIN => \N__50641\,
            DOUT => \N__50640\,
            PACKAGEPIN => test_wire
        );

    \test_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50642\,
            PADOUT => \N__50641\,
            PADIN => \N__50640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50633\,
            DIN => \N__50632\,
            DOUT => \N__50631\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50633\,
            PADOUT => \N__50632\,
            PADIN => \N__50631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50624\,
            DIN => \N__50623\,
            DOUT => \N__50622\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50624\,
            PADOUT => \N__50623\,
            PADIN => \N__50622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50615\,
            DIN => \N__50614\,
            DOUT => \N__50613\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50615\,
            PADOUT => \N__50614\,
            PADIN => \N__50613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50606\,
            DIN => \N__50605\,
            DOUT => \N__50604\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50606\,
            PADOUT => \N__50605\,
            PADIN => \N__50604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50597\,
            DIN => \N__50596\,
            DOUT => \N__50595\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50597\,
            PADOUT => \N__50596\,
            PADIN => \N__50595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test22_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50588\,
            DIN => \N__50587\,
            DOUT => \N__50586\,
            PACKAGEPIN => test22_wire
        );

    \test22_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50588\,
            PADOUT => \N__50587\,
            PADIN => \N__50586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__42400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50579\,
            DIN => \N__50578\,
            DOUT => \N__50577\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50579\,
            PADOUT => \N__50578\,
            PADIN => \N__50577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50570\,
            DIN => \N__50569\,
            DOUT => \N__50568\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50570\,
            PADOUT => \N__50569\,
            PADIN => \N__50568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50561\,
            DIN => \N__50560\,
            DOUT => \N__50559\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50561\,
            PADOUT => \N__50560\,
            PADIN => \N__50559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38920\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50552\,
            DIN => \N__50551\,
            DOUT => \N__50550\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50552\,
            PADOUT => \N__50551\,
            PADIN => \N__50550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50543\,
            DIN => \N__50542\,
            DOUT => \N__50541\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50543\,
            PADOUT => \N__50542\,
            PADIN => \N__50541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28702\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50534\,
            DIN => \N__50533\,
            DOUT => \N__50532\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50534\,
            PADOUT => \N__50533\,
            PADIN => \N__50532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50525\,
            DIN => \N__50524\,
            DOUT => \N__50523\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50525\,
            PADOUT => \N__50524\,
            PADIN => \N__50523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12049\ : CascadeMux
    port map (
            O => \N__50506\,
            I => \N__50502\
        );

    \I__12048\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50498\
        );

    \I__12047\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50495\
        );

    \I__12046\ : InMux
    port map (
            O => \N__50501\,
            I => \N__50492\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__50498\,
            I => \N__50489\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__50495\,
            I => \N__50484\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__50492\,
            I => \N__50484\
        );

    \I__12042\ : Span4Mux_v
    port map (
            O => \N__50489\,
            I => \N__50481\
        );

    \I__12041\ : Span12Mux_v
    port map (
            O => \N__50484\,
            I => \N__50476\
        );

    \I__12040\ : Sp12to4
    port map (
            O => \N__50481\,
            I => \N__50476\
        );

    \I__12039\ : Odrv12
    port map (
            O => \N__50476\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__12038\ : CascadeMux
    port map (
            O => \N__50473\,
            I => \N__50469\
        );

    \I__12037\ : InMux
    port map (
            O => \N__50472\,
            I => \N__50465\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50469\,
            I => \N__50460\
        );

    \I__12035\ : InMux
    port map (
            O => \N__50468\,
            I => \N__50460\
        );

    \I__12034\ : LocalMux
    port map (
            O => \N__50465\,
            I => \N__50457\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__50460\,
            I => pwm_duty_input_7
        );

    \I__12032\ : Odrv4
    port map (
            O => \N__50457\,
            I => pwm_duty_input_7
        );

    \I__12031\ : InMux
    port map (
            O => \N__50452\,
            I => \N__50449\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__50449\,
            I => \N__50446\
        );

    \I__12029\ : Odrv4
    port map (
            O => \N__50446\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50443\,
            I => \N__50434\
        );

    \I__12027\ : InMux
    port map (
            O => \N__50442\,
            I => \N__50434\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50441\,
            I => \N__50434\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__50434\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50431\,
            I => \N__50427\
        );

    \I__12023\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50424\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__50427\,
            I => \N__50421\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__50424\,
            I => pwm_duty_input_0
        );

    \I__12020\ : Odrv4
    port map (
            O => \N__50421\,
            I => pwm_duty_input_0
        );

    \I__12019\ : InMux
    port map (
            O => \N__50416\,
            I => \N__50413\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__50413\,
            I => \N__50409\
        );

    \I__12017\ : InMux
    port map (
            O => \N__50412\,
            I => \N__50406\
        );

    \I__12016\ : Span4Mux_v
    port map (
            O => \N__50409\,
            I => \N__50400\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__50406\,
            I => \N__50400\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50397\
        );

    \I__12013\ : Span4Mux_v
    port map (
            O => \N__50400\,
            I => \N__50394\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50397\,
            I => \N__50391\
        );

    \I__12011\ : Sp12to4
    port map (
            O => \N__50394\,
            I => \N__50388\
        );

    \I__12010\ : Span4Mux_v
    port map (
            O => \N__50391\,
            I => \N__50385\
        );

    \I__12009\ : Span12Mux_s3_h
    port map (
            O => \N__50388\,
            I => \N__50380\
        );

    \I__12008\ : Sp12to4
    port map (
            O => \N__50385\,
            I => \N__50380\
        );

    \I__12007\ : Odrv12
    port map (
            O => \N__50380\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__12006\ : InMux
    port map (
            O => \N__50377\,
            I => \N__50372\
        );

    \I__12005\ : InMux
    port map (
            O => \N__50376\,
            I => \N__50367\
        );

    \I__12004\ : InMux
    port map (
            O => \N__50375\,
            I => \N__50367\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__50372\,
            I => \N__50364\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50367\,
            I => pwm_duty_input_9
        );

    \I__12001\ : Odrv4
    port map (
            O => \N__50364\,
            I => pwm_duty_input_9
        );

    \I__12000\ : CascadeMux
    port map (
            O => \N__50359\,
            I => \N__50356\
        );

    \I__11999\ : InMux
    port map (
            O => \N__50356\,
            I => \N__50353\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50353\,
            I => \N__50349\
        );

    \I__11997\ : InMux
    port map (
            O => \N__50352\,
            I => \N__50346\
        );

    \I__11996\ : Span4Mux_v
    port map (
            O => \N__50349\,
            I => \N__50340\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50346\,
            I => \N__50340\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50345\,
            I => \N__50337\
        );

    \I__11993\ : Span4Mux_v
    port map (
            O => \N__50340\,
            I => \N__50334\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__50337\,
            I => \N__50331\
        );

    \I__11991\ : Sp12to4
    port map (
            O => \N__50334\,
            I => \N__50326\
        );

    \I__11990\ : Span12Mux_v
    port map (
            O => \N__50331\,
            I => \N__50326\
        );

    \I__11989\ : Odrv12
    port map (
            O => \N__50326\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__11988\ : InMux
    port map (
            O => \N__50323\,
            I => \N__50318\
        );

    \I__11987\ : InMux
    port map (
            O => \N__50322\,
            I => \N__50313\
        );

    \I__11986\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50313\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__50318\,
            I => \N__50310\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__50313\,
            I => pwm_duty_input_8
        );

    \I__11983\ : Odrv4
    port map (
            O => \N__50310\,
            I => pwm_duty_input_8
        );

    \I__11982\ : CascadeMux
    port map (
            O => \N__50305\,
            I => \N__50302\
        );

    \I__11981\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50299\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50299\,
            I => \N__50294\
        );

    \I__11979\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50291\
        );

    \I__11978\ : InMux
    port map (
            O => \N__50297\,
            I => \N__50288\
        );

    \I__11977\ : Span4Mux_v
    port map (
            O => \N__50294\,
            I => \N__50283\
        );

    \I__11976\ : LocalMux
    port map (
            O => \N__50291\,
            I => \N__50283\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__50288\,
            I => \N__50280\
        );

    \I__11974\ : Span4Mux_v
    port map (
            O => \N__50283\,
            I => \N__50277\
        );

    \I__11973\ : Span4Mux_v
    port map (
            O => \N__50280\,
            I => \N__50274\
        );

    \I__11972\ : Sp12to4
    port map (
            O => \N__50277\,
            I => \N__50269\
        );

    \I__11971\ : Sp12to4
    port map (
            O => \N__50274\,
            I => \N__50269\
        );

    \I__11970\ : Odrv12
    port map (
            O => \N__50269\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__11969\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50261\
        );

    \I__11968\ : InMux
    port map (
            O => \N__50265\,
            I => \N__50258\
        );

    \I__11967\ : InMux
    port map (
            O => \N__50264\,
            I => \N__50255\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__50261\,
            I => \N__50252\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__50258\,
            I => pwm_duty_input_5
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__50255\,
            I => pwm_duty_input_5
        );

    \I__11963\ : Odrv4
    port map (
            O => \N__50252\,
            I => pwm_duty_input_5
        );

    \I__11962\ : InMux
    port map (
            O => \N__50245\,
            I => \N__50233\
        );

    \I__11961\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50230\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50243\,
            I => \N__50225\
        );

    \I__11959\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50225\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50241\,
            I => \N__50222\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50219\
        );

    \I__11956\ : InMux
    port map (
            O => \N__50239\,
            I => \N__50210\
        );

    \I__11955\ : InMux
    port map (
            O => \N__50238\,
            I => \N__50210\
        );

    \I__11954\ : InMux
    port map (
            O => \N__50237\,
            I => \N__50210\
        );

    \I__11953\ : InMux
    port map (
            O => \N__50236\,
            I => \N__50210\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__50233\,
            I => \N__50203\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__50230\,
            I => \N__50203\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__50225\,
            I => \N__50203\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__50222\,
            I => \N__50200\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__50219\,
            I => \N__50197\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__50210\,
            I => \N__50192\
        );

    \I__11946\ : Sp12to4
    port map (
            O => \N__50203\,
            I => \N__50192\
        );

    \I__11945\ : Span4Mux_h
    port map (
            O => \N__50200\,
            I => \N__50189\
        );

    \I__11944\ : Span12Mux_s1_h
    port map (
            O => \N__50197\,
            I => \N__50184\
        );

    \I__11943\ : Span12Mux_s10_v
    port map (
            O => \N__50192\,
            I => \N__50184\
        );

    \I__11942\ : Odrv4
    port map (
            O => \N__50189\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__11941\ : Odrv12
    port map (
            O => \N__50184\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__11940\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50175\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50171\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__50175\,
            I => \N__50168\
        );

    \I__11937\ : InMux
    port map (
            O => \N__50174\,
            I => \N__50165\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__50171\,
            I => \N__50162\
        );

    \I__11935\ : Span4Mux_v
    port map (
            O => \N__50168\,
            I => \N__50157\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__50165\,
            I => \N__50157\
        );

    \I__11933\ : Span4Mux_v
    port map (
            O => \N__50162\,
            I => \N__50154\
        );

    \I__11932\ : Span4Mux_v
    port map (
            O => \N__50157\,
            I => \N__50151\
        );

    \I__11931\ : Sp12to4
    port map (
            O => \N__50154\,
            I => \N__50146\
        );

    \I__11930\ : Sp12to4
    port map (
            O => \N__50151\,
            I => \N__50146\
        );

    \I__11929\ : Odrv12
    port map (
            O => \N__50146\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__11928\ : CascadeMux
    port map (
            O => \N__50143\,
            I => \N__50137\
        );

    \I__11927\ : CascadeMux
    port map (
            O => \N__50142\,
            I => \N__50134\
        );

    \I__11926\ : InMux
    port map (
            O => \N__50141\,
            I => \N__50125\
        );

    \I__11925\ : InMux
    port map (
            O => \N__50140\,
            I => \N__50125\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50125\
        );

    \I__11923\ : InMux
    port map (
            O => \N__50134\,
            I => \N__50125\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__50125\,
            I => \N__50118\
        );

    \I__11921\ : InMux
    port map (
            O => \N__50124\,
            I => \N__50115\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50123\,
            I => \N__50110\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50122\,
            I => \N__50110\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50121\,
            I => \N__50107\
        );

    \I__11917\ : Span4Mux_s2_h
    port map (
            O => \N__50118\,
            I => \N__50100\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__50115\,
            I => \N__50100\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__50110\,
            I => \N__50100\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__50107\,
            I => \N__50097\
        );

    \I__11913\ : Span4Mux_v
    port map (
            O => \N__50100\,
            I => \N__50094\
        );

    \I__11912\ : Span12Mux_s10_h
    port map (
            O => \N__50097\,
            I => \N__50091\
        );

    \I__11911\ : Span4Mux_h
    port map (
            O => \N__50094\,
            I => \N__50088\
        );

    \I__11910\ : Odrv12
    port map (
            O => \N__50091\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__11909\ : Odrv4
    port map (
            O => \N__50088\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__11908\ : InMux
    port map (
            O => \N__50083\,
            I => \N__50069\
        );

    \I__11907\ : InMux
    port map (
            O => \N__50082\,
            I => \N__50069\
        );

    \I__11906\ : InMux
    port map (
            O => \N__50081\,
            I => \N__50069\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50080\,
            I => \N__50069\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50079\,
            I => \N__50064\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50078\,
            I => \N__50064\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__50069\,
            I => \N__50058\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__50064\,
            I => \N__50058\
        );

    \I__11900\ : InMux
    port map (
            O => \N__50063\,
            I => \N__50055\
        );

    \I__11899\ : Span4Mux_v
    port map (
            O => \N__50058\,
            I => \N__50050\
        );

    \I__11898\ : LocalMux
    port map (
            O => \N__50055\,
            I => \N__50050\
        );

    \I__11897\ : Span4Mux_h
    port map (
            O => \N__50050\,
            I => \N__50047\
        );

    \I__11896\ : Span4Mux_h
    port map (
            O => \N__50047\,
            I => \N__50044\
        );

    \I__11895\ : Odrv4
    port map (
            O => \N__50044\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__11894\ : InMux
    port map (
            O => \N__50041\,
            I => \N__50036\
        );

    \I__11893\ : InMux
    port map (
            O => \N__50040\,
            I => \N__50031\
        );

    \I__11892\ : InMux
    port map (
            O => \N__50039\,
            I => \N__50031\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__50036\,
            I => \N__50028\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__50031\,
            I => pwm_duty_input_6
        );

    \I__11889\ : Odrv4
    port map (
            O => \N__50028\,
            I => pwm_duty_input_6
        );

    \I__11888\ : InMux
    port map (
            O => \N__50023\,
            I => \N__50020\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__50020\,
            I => \N__49869\
        );

    \I__11886\ : ClkMux
    port map (
            O => \N__50019\,
            I => \N__49558\
        );

    \I__11885\ : ClkMux
    port map (
            O => \N__50018\,
            I => \N__49558\
        );

    \I__11884\ : ClkMux
    port map (
            O => \N__50017\,
            I => \N__49558\
        );

    \I__11883\ : ClkMux
    port map (
            O => \N__50016\,
            I => \N__49558\
        );

    \I__11882\ : ClkMux
    port map (
            O => \N__50015\,
            I => \N__49558\
        );

    \I__11881\ : ClkMux
    port map (
            O => \N__50014\,
            I => \N__49558\
        );

    \I__11880\ : ClkMux
    port map (
            O => \N__50013\,
            I => \N__49558\
        );

    \I__11879\ : ClkMux
    port map (
            O => \N__50012\,
            I => \N__49558\
        );

    \I__11878\ : ClkMux
    port map (
            O => \N__50011\,
            I => \N__49558\
        );

    \I__11877\ : ClkMux
    port map (
            O => \N__50010\,
            I => \N__49558\
        );

    \I__11876\ : ClkMux
    port map (
            O => \N__50009\,
            I => \N__49558\
        );

    \I__11875\ : ClkMux
    port map (
            O => \N__50008\,
            I => \N__49558\
        );

    \I__11874\ : ClkMux
    port map (
            O => \N__50007\,
            I => \N__49558\
        );

    \I__11873\ : ClkMux
    port map (
            O => \N__50006\,
            I => \N__49558\
        );

    \I__11872\ : ClkMux
    port map (
            O => \N__50005\,
            I => \N__49558\
        );

    \I__11871\ : ClkMux
    port map (
            O => \N__50004\,
            I => \N__49558\
        );

    \I__11870\ : ClkMux
    port map (
            O => \N__50003\,
            I => \N__49558\
        );

    \I__11869\ : ClkMux
    port map (
            O => \N__50002\,
            I => \N__49558\
        );

    \I__11868\ : ClkMux
    port map (
            O => \N__50001\,
            I => \N__49558\
        );

    \I__11867\ : ClkMux
    port map (
            O => \N__50000\,
            I => \N__49558\
        );

    \I__11866\ : ClkMux
    port map (
            O => \N__49999\,
            I => \N__49558\
        );

    \I__11865\ : ClkMux
    port map (
            O => \N__49998\,
            I => \N__49558\
        );

    \I__11864\ : ClkMux
    port map (
            O => \N__49997\,
            I => \N__49558\
        );

    \I__11863\ : ClkMux
    port map (
            O => \N__49996\,
            I => \N__49558\
        );

    \I__11862\ : ClkMux
    port map (
            O => \N__49995\,
            I => \N__49558\
        );

    \I__11861\ : ClkMux
    port map (
            O => \N__49994\,
            I => \N__49558\
        );

    \I__11860\ : ClkMux
    port map (
            O => \N__49993\,
            I => \N__49558\
        );

    \I__11859\ : ClkMux
    port map (
            O => \N__49992\,
            I => \N__49558\
        );

    \I__11858\ : ClkMux
    port map (
            O => \N__49991\,
            I => \N__49558\
        );

    \I__11857\ : ClkMux
    port map (
            O => \N__49990\,
            I => \N__49558\
        );

    \I__11856\ : ClkMux
    port map (
            O => \N__49989\,
            I => \N__49558\
        );

    \I__11855\ : ClkMux
    port map (
            O => \N__49988\,
            I => \N__49558\
        );

    \I__11854\ : ClkMux
    port map (
            O => \N__49987\,
            I => \N__49558\
        );

    \I__11853\ : ClkMux
    port map (
            O => \N__49986\,
            I => \N__49558\
        );

    \I__11852\ : ClkMux
    port map (
            O => \N__49985\,
            I => \N__49558\
        );

    \I__11851\ : ClkMux
    port map (
            O => \N__49984\,
            I => \N__49558\
        );

    \I__11850\ : ClkMux
    port map (
            O => \N__49983\,
            I => \N__49558\
        );

    \I__11849\ : ClkMux
    port map (
            O => \N__49982\,
            I => \N__49558\
        );

    \I__11848\ : ClkMux
    port map (
            O => \N__49981\,
            I => \N__49558\
        );

    \I__11847\ : ClkMux
    port map (
            O => \N__49980\,
            I => \N__49558\
        );

    \I__11846\ : ClkMux
    port map (
            O => \N__49979\,
            I => \N__49558\
        );

    \I__11845\ : ClkMux
    port map (
            O => \N__49978\,
            I => \N__49558\
        );

    \I__11844\ : ClkMux
    port map (
            O => \N__49977\,
            I => \N__49558\
        );

    \I__11843\ : ClkMux
    port map (
            O => \N__49976\,
            I => \N__49558\
        );

    \I__11842\ : ClkMux
    port map (
            O => \N__49975\,
            I => \N__49558\
        );

    \I__11841\ : ClkMux
    port map (
            O => \N__49974\,
            I => \N__49558\
        );

    \I__11840\ : ClkMux
    port map (
            O => \N__49973\,
            I => \N__49558\
        );

    \I__11839\ : ClkMux
    port map (
            O => \N__49972\,
            I => \N__49558\
        );

    \I__11838\ : ClkMux
    port map (
            O => \N__49971\,
            I => \N__49558\
        );

    \I__11837\ : ClkMux
    port map (
            O => \N__49970\,
            I => \N__49558\
        );

    \I__11836\ : ClkMux
    port map (
            O => \N__49969\,
            I => \N__49558\
        );

    \I__11835\ : ClkMux
    port map (
            O => \N__49968\,
            I => \N__49558\
        );

    \I__11834\ : ClkMux
    port map (
            O => \N__49967\,
            I => \N__49558\
        );

    \I__11833\ : ClkMux
    port map (
            O => \N__49966\,
            I => \N__49558\
        );

    \I__11832\ : ClkMux
    port map (
            O => \N__49965\,
            I => \N__49558\
        );

    \I__11831\ : ClkMux
    port map (
            O => \N__49964\,
            I => \N__49558\
        );

    \I__11830\ : ClkMux
    port map (
            O => \N__49963\,
            I => \N__49558\
        );

    \I__11829\ : ClkMux
    port map (
            O => \N__49962\,
            I => \N__49558\
        );

    \I__11828\ : ClkMux
    port map (
            O => \N__49961\,
            I => \N__49558\
        );

    \I__11827\ : ClkMux
    port map (
            O => \N__49960\,
            I => \N__49558\
        );

    \I__11826\ : ClkMux
    port map (
            O => \N__49959\,
            I => \N__49558\
        );

    \I__11825\ : ClkMux
    port map (
            O => \N__49958\,
            I => \N__49558\
        );

    \I__11824\ : ClkMux
    port map (
            O => \N__49957\,
            I => \N__49558\
        );

    \I__11823\ : ClkMux
    port map (
            O => \N__49956\,
            I => \N__49558\
        );

    \I__11822\ : ClkMux
    port map (
            O => \N__49955\,
            I => \N__49558\
        );

    \I__11821\ : ClkMux
    port map (
            O => \N__49954\,
            I => \N__49558\
        );

    \I__11820\ : ClkMux
    port map (
            O => \N__49953\,
            I => \N__49558\
        );

    \I__11819\ : ClkMux
    port map (
            O => \N__49952\,
            I => \N__49558\
        );

    \I__11818\ : ClkMux
    port map (
            O => \N__49951\,
            I => \N__49558\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__49950\,
            I => \N__49558\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__49949\,
            I => \N__49558\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__49948\,
            I => \N__49558\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__49947\,
            I => \N__49558\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__49946\,
            I => \N__49558\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__49945\,
            I => \N__49558\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__49944\,
            I => \N__49558\
        );

    \I__11810\ : ClkMux
    port map (
            O => \N__49943\,
            I => \N__49558\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__49942\,
            I => \N__49558\
        );

    \I__11808\ : ClkMux
    port map (
            O => \N__49941\,
            I => \N__49558\
        );

    \I__11807\ : ClkMux
    port map (
            O => \N__49940\,
            I => \N__49558\
        );

    \I__11806\ : ClkMux
    port map (
            O => \N__49939\,
            I => \N__49558\
        );

    \I__11805\ : ClkMux
    port map (
            O => \N__49938\,
            I => \N__49558\
        );

    \I__11804\ : ClkMux
    port map (
            O => \N__49937\,
            I => \N__49558\
        );

    \I__11803\ : ClkMux
    port map (
            O => \N__49936\,
            I => \N__49558\
        );

    \I__11802\ : ClkMux
    port map (
            O => \N__49935\,
            I => \N__49558\
        );

    \I__11801\ : ClkMux
    port map (
            O => \N__49934\,
            I => \N__49558\
        );

    \I__11800\ : ClkMux
    port map (
            O => \N__49933\,
            I => \N__49558\
        );

    \I__11799\ : ClkMux
    port map (
            O => \N__49932\,
            I => \N__49558\
        );

    \I__11798\ : ClkMux
    port map (
            O => \N__49931\,
            I => \N__49558\
        );

    \I__11797\ : ClkMux
    port map (
            O => \N__49930\,
            I => \N__49558\
        );

    \I__11796\ : ClkMux
    port map (
            O => \N__49929\,
            I => \N__49558\
        );

    \I__11795\ : ClkMux
    port map (
            O => \N__49928\,
            I => \N__49558\
        );

    \I__11794\ : ClkMux
    port map (
            O => \N__49927\,
            I => \N__49558\
        );

    \I__11793\ : ClkMux
    port map (
            O => \N__49926\,
            I => \N__49558\
        );

    \I__11792\ : ClkMux
    port map (
            O => \N__49925\,
            I => \N__49558\
        );

    \I__11791\ : ClkMux
    port map (
            O => \N__49924\,
            I => \N__49558\
        );

    \I__11790\ : ClkMux
    port map (
            O => \N__49923\,
            I => \N__49558\
        );

    \I__11789\ : ClkMux
    port map (
            O => \N__49922\,
            I => \N__49558\
        );

    \I__11788\ : ClkMux
    port map (
            O => \N__49921\,
            I => \N__49558\
        );

    \I__11787\ : ClkMux
    port map (
            O => \N__49920\,
            I => \N__49558\
        );

    \I__11786\ : ClkMux
    port map (
            O => \N__49919\,
            I => \N__49558\
        );

    \I__11785\ : ClkMux
    port map (
            O => \N__49918\,
            I => \N__49558\
        );

    \I__11784\ : ClkMux
    port map (
            O => \N__49917\,
            I => \N__49558\
        );

    \I__11783\ : ClkMux
    port map (
            O => \N__49916\,
            I => \N__49558\
        );

    \I__11782\ : ClkMux
    port map (
            O => \N__49915\,
            I => \N__49558\
        );

    \I__11781\ : ClkMux
    port map (
            O => \N__49914\,
            I => \N__49558\
        );

    \I__11780\ : ClkMux
    port map (
            O => \N__49913\,
            I => \N__49558\
        );

    \I__11779\ : ClkMux
    port map (
            O => \N__49912\,
            I => \N__49558\
        );

    \I__11778\ : ClkMux
    port map (
            O => \N__49911\,
            I => \N__49558\
        );

    \I__11777\ : ClkMux
    port map (
            O => \N__49910\,
            I => \N__49558\
        );

    \I__11776\ : ClkMux
    port map (
            O => \N__49909\,
            I => \N__49558\
        );

    \I__11775\ : ClkMux
    port map (
            O => \N__49908\,
            I => \N__49558\
        );

    \I__11774\ : ClkMux
    port map (
            O => \N__49907\,
            I => \N__49558\
        );

    \I__11773\ : ClkMux
    port map (
            O => \N__49906\,
            I => \N__49558\
        );

    \I__11772\ : ClkMux
    port map (
            O => \N__49905\,
            I => \N__49558\
        );

    \I__11771\ : ClkMux
    port map (
            O => \N__49904\,
            I => \N__49558\
        );

    \I__11770\ : ClkMux
    port map (
            O => \N__49903\,
            I => \N__49558\
        );

    \I__11769\ : ClkMux
    port map (
            O => \N__49902\,
            I => \N__49558\
        );

    \I__11768\ : ClkMux
    port map (
            O => \N__49901\,
            I => \N__49558\
        );

    \I__11767\ : ClkMux
    port map (
            O => \N__49900\,
            I => \N__49558\
        );

    \I__11766\ : ClkMux
    port map (
            O => \N__49899\,
            I => \N__49558\
        );

    \I__11765\ : ClkMux
    port map (
            O => \N__49898\,
            I => \N__49558\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__49897\,
            I => \N__49558\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__49896\,
            I => \N__49558\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__49895\,
            I => \N__49558\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__49894\,
            I => \N__49558\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__49893\,
            I => \N__49558\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__49892\,
            I => \N__49558\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__49891\,
            I => \N__49558\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__49890\,
            I => \N__49558\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__49889\,
            I => \N__49558\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__49888\,
            I => \N__49558\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__49887\,
            I => \N__49558\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__49886\,
            I => \N__49558\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__49885\,
            I => \N__49558\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__49884\,
            I => \N__49558\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__49883\,
            I => \N__49558\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__49882\,
            I => \N__49558\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__49881\,
            I => \N__49558\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__49880\,
            I => \N__49558\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__49879\,
            I => \N__49558\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__49878\,
            I => \N__49558\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__49877\,
            I => \N__49558\
        );

    \I__11743\ : ClkMux
    port map (
            O => \N__49876\,
            I => \N__49558\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__49875\,
            I => \N__49558\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__49874\,
            I => \N__49558\
        );

    \I__11740\ : ClkMux
    port map (
            O => \N__49873\,
            I => \N__49558\
        );

    \I__11739\ : ClkMux
    port map (
            O => \N__49872\,
            I => \N__49558\
        );

    \I__11738\ : Glb2LocalMux
    port map (
            O => \N__49869\,
            I => \N__49558\
        );

    \I__11737\ : ClkMux
    port map (
            O => \N__49868\,
            I => \N__49558\
        );

    \I__11736\ : ClkMux
    port map (
            O => \N__49867\,
            I => \N__49558\
        );

    \I__11735\ : ClkMux
    port map (
            O => \N__49866\,
            I => \N__49558\
        );

    \I__11734\ : ClkMux
    port map (
            O => \N__49865\,
            I => \N__49558\
        );

    \I__11733\ : GlobalMux
    port map (
            O => \N__49558\,
            I => clock_output_0
        );

    \I__11732\ : InMux
    port map (
            O => \N__49555\,
            I => \N__49549\
        );

    \I__11731\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49546\
        );

    \I__11730\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49543\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49552\,
            I => \N__49540\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__49549\,
            I => \N__49537\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49534\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__49543\,
            I => \N__49531\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__49540\,
            I => \N__49527\
        );

    \I__11724\ : Glb2LocalMux
    port map (
            O => \N__49537\,
            I => \N__49057\
        );

    \I__11723\ : Glb2LocalMux
    port map (
            O => \N__49534\,
            I => \N__49057\
        );

    \I__11722\ : Glb2LocalMux
    port map (
            O => \N__49531\,
            I => \N__49057\
        );

    \I__11721\ : SRMux
    port map (
            O => \N__49530\,
            I => \N__49057\
        );

    \I__11720\ : Glb2LocalMux
    port map (
            O => \N__49527\,
            I => \N__49057\
        );

    \I__11719\ : SRMux
    port map (
            O => \N__49526\,
            I => \N__49057\
        );

    \I__11718\ : SRMux
    port map (
            O => \N__49525\,
            I => \N__49057\
        );

    \I__11717\ : SRMux
    port map (
            O => \N__49524\,
            I => \N__49057\
        );

    \I__11716\ : SRMux
    port map (
            O => \N__49523\,
            I => \N__49057\
        );

    \I__11715\ : SRMux
    port map (
            O => \N__49522\,
            I => \N__49057\
        );

    \I__11714\ : SRMux
    port map (
            O => \N__49521\,
            I => \N__49057\
        );

    \I__11713\ : SRMux
    port map (
            O => \N__49520\,
            I => \N__49057\
        );

    \I__11712\ : SRMux
    port map (
            O => \N__49519\,
            I => \N__49057\
        );

    \I__11711\ : SRMux
    port map (
            O => \N__49518\,
            I => \N__49057\
        );

    \I__11710\ : SRMux
    port map (
            O => \N__49517\,
            I => \N__49057\
        );

    \I__11709\ : SRMux
    port map (
            O => \N__49516\,
            I => \N__49057\
        );

    \I__11708\ : SRMux
    port map (
            O => \N__49515\,
            I => \N__49057\
        );

    \I__11707\ : SRMux
    port map (
            O => \N__49514\,
            I => \N__49057\
        );

    \I__11706\ : SRMux
    port map (
            O => \N__49513\,
            I => \N__49057\
        );

    \I__11705\ : SRMux
    port map (
            O => \N__49512\,
            I => \N__49057\
        );

    \I__11704\ : SRMux
    port map (
            O => \N__49511\,
            I => \N__49057\
        );

    \I__11703\ : SRMux
    port map (
            O => \N__49510\,
            I => \N__49057\
        );

    \I__11702\ : SRMux
    port map (
            O => \N__49509\,
            I => \N__49057\
        );

    \I__11701\ : SRMux
    port map (
            O => \N__49508\,
            I => \N__49057\
        );

    \I__11700\ : SRMux
    port map (
            O => \N__49507\,
            I => \N__49057\
        );

    \I__11699\ : SRMux
    port map (
            O => \N__49506\,
            I => \N__49057\
        );

    \I__11698\ : SRMux
    port map (
            O => \N__49505\,
            I => \N__49057\
        );

    \I__11697\ : SRMux
    port map (
            O => \N__49504\,
            I => \N__49057\
        );

    \I__11696\ : SRMux
    port map (
            O => \N__49503\,
            I => \N__49057\
        );

    \I__11695\ : SRMux
    port map (
            O => \N__49502\,
            I => \N__49057\
        );

    \I__11694\ : SRMux
    port map (
            O => \N__49501\,
            I => \N__49057\
        );

    \I__11693\ : SRMux
    port map (
            O => \N__49500\,
            I => \N__49057\
        );

    \I__11692\ : SRMux
    port map (
            O => \N__49499\,
            I => \N__49057\
        );

    \I__11691\ : SRMux
    port map (
            O => \N__49498\,
            I => \N__49057\
        );

    \I__11690\ : SRMux
    port map (
            O => \N__49497\,
            I => \N__49057\
        );

    \I__11689\ : SRMux
    port map (
            O => \N__49496\,
            I => \N__49057\
        );

    \I__11688\ : SRMux
    port map (
            O => \N__49495\,
            I => \N__49057\
        );

    \I__11687\ : SRMux
    port map (
            O => \N__49494\,
            I => \N__49057\
        );

    \I__11686\ : SRMux
    port map (
            O => \N__49493\,
            I => \N__49057\
        );

    \I__11685\ : SRMux
    port map (
            O => \N__49492\,
            I => \N__49057\
        );

    \I__11684\ : SRMux
    port map (
            O => \N__49491\,
            I => \N__49057\
        );

    \I__11683\ : SRMux
    port map (
            O => \N__49490\,
            I => \N__49057\
        );

    \I__11682\ : SRMux
    port map (
            O => \N__49489\,
            I => \N__49057\
        );

    \I__11681\ : SRMux
    port map (
            O => \N__49488\,
            I => \N__49057\
        );

    \I__11680\ : SRMux
    port map (
            O => \N__49487\,
            I => \N__49057\
        );

    \I__11679\ : SRMux
    port map (
            O => \N__49486\,
            I => \N__49057\
        );

    \I__11678\ : SRMux
    port map (
            O => \N__49485\,
            I => \N__49057\
        );

    \I__11677\ : SRMux
    port map (
            O => \N__49484\,
            I => \N__49057\
        );

    \I__11676\ : SRMux
    port map (
            O => \N__49483\,
            I => \N__49057\
        );

    \I__11675\ : SRMux
    port map (
            O => \N__49482\,
            I => \N__49057\
        );

    \I__11674\ : SRMux
    port map (
            O => \N__49481\,
            I => \N__49057\
        );

    \I__11673\ : SRMux
    port map (
            O => \N__49480\,
            I => \N__49057\
        );

    \I__11672\ : SRMux
    port map (
            O => \N__49479\,
            I => \N__49057\
        );

    \I__11671\ : SRMux
    port map (
            O => \N__49478\,
            I => \N__49057\
        );

    \I__11670\ : SRMux
    port map (
            O => \N__49477\,
            I => \N__49057\
        );

    \I__11669\ : SRMux
    port map (
            O => \N__49476\,
            I => \N__49057\
        );

    \I__11668\ : SRMux
    port map (
            O => \N__49475\,
            I => \N__49057\
        );

    \I__11667\ : SRMux
    port map (
            O => \N__49474\,
            I => \N__49057\
        );

    \I__11666\ : SRMux
    port map (
            O => \N__49473\,
            I => \N__49057\
        );

    \I__11665\ : SRMux
    port map (
            O => \N__49472\,
            I => \N__49057\
        );

    \I__11664\ : SRMux
    port map (
            O => \N__49471\,
            I => \N__49057\
        );

    \I__11663\ : SRMux
    port map (
            O => \N__49470\,
            I => \N__49057\
        );

    \I__11662\ : SRMux
    port map (
            O => \N__49469\,
            I => \N__49057\
        );

    \I__11661\ : SRMux
    port map (
            O => \N__49468\,
            I => \N__49057\
        );

    \I__11660\ : SRMux
    port map (
            O => \N__49467\,
            I => \N__49057\
        );

    \I__11659\ : SRMux
    port map (
            O => \N__49466\,
            I => \N__49057\
        );

    \I__11658\ : SRMux
    port map (
            O => \N__49465\,
            I => \N__49057\
        );

    \I__11657\ : SRMux
    port map (
            O => \N__49464\,
            I => \N__49057\
        );

    \I__11656\ : SRMux
    port map (
            O => \N__49463\,
            I => \N__49057\
        );

    \I__11655\ : SRMux
    port map (
            O => \N__49462\,
            I => \N__49057\
        );

    \I__11654\ : SRMux
    port map (
            O => \N__49461\,
            I => \N__49057\
        );

    \I__11653\ : SRMux
    port map (
            O => \N__49460\,
            I => \N__49057\
        );

    \I__11652\ : SRMux
    port map (
            O => \N__49459\,
            I => \N__49057\
        );

    \I__11651\ : SRMux
    port map (
            O => \N__49458\,
            I => \N__49057\
        );

    \I__11650\ : SRMux
    port map (
            O => \N__49457\,
            I => \N__49057\
        );

    \I__11649\ : SRMux
    port map (
            O => \N__49456\,
            I => \N__49057\
        );

    \I__11648\ : SRMux
    port map (
            O => \N__49455\,
            I => \N__49057\
        );

    \I__11647\ : SRMux
    port map (
            O => \N__49454\,
            I => \N__49057\
        );

    \I__11646\ : SRMux
    port map (
            O => \N__49453\,
            I => \N__49057\
        );

    \I__11645\ : SRMux
    port map (
            O => \N__49452\,
            I => \N__49057\
        );

    \I__11644\ : SRMux
    port map (
            O => \N__49451\,
            I => \N__49057\
        );

    \I__11643\ : SRMux
    port map (
            O => \N__49450\,
            I => \N__49057\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__49449\,
            I => \N__49057\
        );

    \I__11641\ : SRMux
    port map (
            O => \N__49448\,
            I => \N__49057\
        );

    \I__11640\ : SRMux
    port map (
            O => \N__49447\,
            I => \N__49057\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__49446\,
            I => \N__49057\
        );

    \I__11638\ : SRMux
    port map (
            O => \N__49445\,
            I => \N__49057\
        );

    \I__11637\ : SRMux
    port map (
            O => \N__49444\,
            I => \N__49057\
        );

    \I__11636\ : SRMux
    port map (
            O => \N__49443\,
            I => \N__49057\
        );

    \I__11635\ : SRMux
    port map (
            O => \N__49442\,
            I => \N__49057\
        );

    \I__11634\ : SRMux
    port map (
            O => \N__49441\,
            I => \N__49057\
        );

    \I__11633\ : SRMux
    port map (
            O => \N__49440\,
            I => \N__49057\
        );

    \I__11632\ : SRMux
    port map (
            O => \N__49439\,
            I => \N__49057\
        );

    \I__11631\ : SRMux
    port map (
            O => \N__49438\,
            I => \N__49057\
        );

    \I__11630\ : SRMux
    port map (
            O => \N__49437\,
            I => \N__49057\
        );

    \I__11629\ : SRMux
    port map (
            O => \N__49436\,
            I => \N__49057\
        );

    \I__11628\ : SRMux
    port map (
            O => \N__49435\,
            I => \N__49057\
        );

    \I__11627\ : SRMux
    port map (
            O => \N__49434\,
            I => \N__49057\
        );

    \I__11626\ : SRMux
    port map (
            O => \N__49433\,
            I => \N__49057\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49432\,
            I => \N__49057\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49431\,
            I => \N__49057\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49430\,
            I => \N__49057\
        );

    \I__11622\ : SRMux
    port map (
            O => \N__49429\,
            I => \N__49057\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49428\,
            I => \N__49057\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49427\,
            I => \N__49057\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49426\,
            I => \N__49057\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49425\,
            I => \N__49057\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49424\,
            I => \N__49057\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49423\,
            I => \N__49057\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49422\,
            I => \N__49057\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49421\,
            I => \N__49057\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49420\,
            I => \N__49057\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49419\,
            I => \N__49057\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49418\,
            I => \N__49057\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49417\,
            I => \N__49057\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49416\,
            I => \N__49057\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49415\,
            I => \N__49057\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49414\,
            I => \N__49057\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49413\,
            I => \N__49057\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49412\,
            I => \N__49057\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49411\,
            I => \N__49057\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49410\,
            I => \N__49057\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49409\,
            I => \N__49057\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49408\,
            I => \N__49057\
        );

    \I__11600\ : SRMux
    port map (
            O => \N__49407\,
            I => \N__49057\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49406\,
            I => \N__49057\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49405\,
            I => \N__49057\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49404\,
            I => \N__49057\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49403\,
            I => \N__49057\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49402\,
            I => \N__49057\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49401\,
            I => \N__49057\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49400\,
            I => \N__49057\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49399\,
            I => \N__49057\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49398\,
            I => \N__49057\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49397\,
            I => \N__49057\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49396\,
            I => \N__49057\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49395\,
            I => \N__49057\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49394\,
            I => \N__49057\
        );

    \I__11586\ : SRMux
    port map (
            O => \N__49393\,
            I => \N__49057\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49392\,
            I => \N__49057\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49391\,
            I => \N__49057\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49390\,
            I => \N__49057\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49389\,
            I => \N__49057\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49388\,
            I => \N__49057\
        );

    \I__11580\ : SRMux
    port map (
            O => \N__49387\,
            I => \N__49057\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49386\,
            I => \N__49057\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49385\,
            I => \N__49057\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49384\,
            I => \N__49057\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49383\,
            I => \N__49057\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49382\,
            I => \N__49057\
        );

    \I__11574\ : SRMux
    port map (
            O => \N__49381\,
            I => \N__49057\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49380\,
            I => \N__49057\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49379\,
            I => \N__49057\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49378\,
            I => \N__49057\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49377\,
            I => \N__49057\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49376\,
            I => \N__49057\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49375\,
            I => \N__49057\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49374\,
            I => \N__49057\
        );

    \I__11566\ : GlobalMux
    port map (
            O => \N__49057\,
            I => \N__49054\
        );

    \I__11565\ : gio2CtrlBuf
    port map (
            O => \N__49054\,
            I => red_c_g
        );

    \I__11564\ : InMux
    port map (
            O => \N__49051\,
            I => \N__49048\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__49048\,
            I => \N__49038\
        );

    \I__11562\ : InMux
    port map (
            O => \N__49047\,
            I => \N__49023\
        );

    \I__11561\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49023\
        );

    \I__11560\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49023\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49023\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49043\,
            I => \N__49023\
        );

    \I__11557\ : InMux
    port map (
            O => \N__49042\,
            I => \N__49023\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49041\,
            I => \N__49023\
        );

    \I__11555\ : Span4Mux_v
    port map (
            O => \N__49038\,
            I => \N__49018\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__49023\,
            I => \N__49018\
        );

    \I__11553\ : Span4Mux_v
    port map (
            O => \N__49018\,
            I => \N__49013\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49017\,
            I => \N__49008\
        );

    \I__11551\ : InMux
    port map (
            O => \N__49016\,
            I => \N__49008\
        );

    \I__11550\ : Sp12to4
    port map (
            O => \N__49013\,
            I => \N__49003\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__49003\
        );

    \I__11548\ : Span12Mux_h
    port map (
            O => \N__49003\,
            I => \N__49000\
        );

    \I__11547\ : Odrv12
    port map (
            O => \N__49000\,
            I => \pwm_generator_inst.N_17\
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__48997\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__11545\ : InMux
    port map (
            O => \N__48994\,
            I => \N__48991\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__48991\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__11543\ : CascadeMux
    port map (
            O => \N__48988\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \I__11542\ : CascadeMux
    port map (
            O => \N__48985\,
            I => \N__48982\
        );

    \I__11541\ : InMux
    port map (
            O => \N__48982\,
            I => \N__48979\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__48979\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__11539\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48973\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__48973\,
            I => \N__48970\
        );

    \I__11537\ : Span4Mux_v
    port map (
            O => \N__48970\,
            I => \N__48967\
        );

    \I__11536\ : Sp12to4
    port map (
            O => \N__48967\,
            I => \N__48964\
        );

    \I__11535\ : Span12Mux_s11_h
    port map (
            O => \N__48964\,
            I => \N__48961\
        );

    \I__11534\ : Odrv12
    port map (
            O => \N__48961\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__11533\ : InMux
    port map (
            O => \N__48958\,
            I => \N__48955\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__48955\,
            I => \N__48951\
        );

    \I__11531\ : InMux
    port map (
            O => \N__48954\,
            I => \N__48948\
        );

    \I__11530\ : Span4Mux_v
    port map (
            O => \N__48951\,
            I => \N__48945\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__48948\,
            I => pwm_duty_input_2
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__48945\,
            I => pwm_duty_input_2
        );

    \I__11527\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48937\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48934\
        );

    \I__11525\ : Odrv4
    port map (
            O => \N__48934\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__11524\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48928\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__48928\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__11522\ : CascadeMux
    port map (
            O => \N__48925\,
            I => \N__48920\
        );

    \I__11521\ : CascadeMux
    port map (
            O => \N__48924\,
            I => \N__48917\
        );

    \I__11520\ : CascadeMux
    port map (
            O => \N__48923\,
            I => \N__48914\
        );

    \I__11519\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48911\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48917\,
            I => \N__48908\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48914\,
            I => \N__48905\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__48911\,
            I => \N__48898\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__48908\,
            I => \N__48898\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__48905\,
            I => \N__48898\
        );

    \I__11513\ : Span4Mux_v
    port map (
            O => \N__48898\,
            I => \N__48894\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48897\,
            I => \N__48891\
        );

    \I__11511\ : Sp12to4
    port map (
            O => \N__48894\,
            I => \N__48886\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__48891\,
            I => \N__48886\
        );

    \I__11509\ : Span12Mux_s11_h
    port map (
            O => \N__48886\,
            I => \N__48883\
        );

    \I__11508\ : Odrv12
    port map (
            O => \N__48883\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__11507\ : CascadeMux
    port map (
            O => \N__48880\,
            I => \N__48877\
        );

    \I__11506\ : InMux
    port map (
            O => \N__48877\,
            I => \N__48872\
        );

    \I__11505\ : CascadeMux
    port map (
            O => \N__48876\,
            I => \N__48869\
        );

    \I__11504\ : InMux
    port map (
            O => \N__48875\,
            I => \N__48866\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__48872\,
            I => \N__48863\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48860\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48866\,
            I => \N__48857\
        );

    \I__11500\ : Span4Mux_h
    port map (
            O => \N__48863\,
            I => \N__48854\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__48860\,
            I => \N__48851\
        );

    \I__11498\ : Span4Mux_v
    port map (
            O => \N__48857\,
            I => \N__48848\
        );

    \I__11497\ : Odrv4
    port map (
            O => \N__48854\,
            I => pwm_duty_input_4
        );

    \I__11496\ : Odrv4
    port map (
            O => \N__48851\,
            I => pwm_duty_input_4
        );

    \I__11495\ : Odrv4
    port map (
            O => \N__48848\,
            I => pwm_duty_input_4
        );

    \I__11494\ : InMux
    port map (
            O => \N__48841\,
            I => \N__48838\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__48838\,
            I => \N__48835\
        );

    \I__11492\ : Span4Mux_v
    port map (
            O => \N__48835\,
            I => \N__48832\
        );

    \I__11491\ : Span4Mux_h
    port map (
            O => \N__48832\,
            I => \N__48829\
        );

    \I__11490\ : Span4Mux_h
    port map (
            O => \N__48829\,
            I => \N__48826\
        );

    \I__11489\ : Odrv4
    port map (
            O => \N__48826\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48823\,
            I => \N__48820\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__48820\,
            I => \N__48816\
        );

    \I__11486\ : InMux
    port map (
            O => \N__48819\,
            I => \N__48813\
        );

    \I__11485\ : Span4Mux_s1_h
    port map (
            O => \N__48816\,
            I => \N__48810\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__48813\,
            I => pwm_duty_input_1
        );

    \I__11483\ : Odrv4
    port map (
            O => \N__48810\,
            I => pwm_duty_input_1
        );

    \I__11482\ : InMux
    port map (
            O => \N__48805\,
            I => \N__48802\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__48802\,
            I => \N__48799\
        );

    \I__11480\ : Span4Mux_v
    port map (
            O => \N__48799\,
            I => \N__48795\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48792\
        );

    \I__11478\ : Odrv4
    port map (
            O => \N__48795\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48792\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48783\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48786\,
            I => \N__48780\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__48783\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__48780\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48770\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48767\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48773\,
            I => \N__48764\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48761\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__48767\,
            I => \N__48758\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48755\
        );

    \I__11466\ : Span4Mux_v
    port map (
            O => \N__48761\,
            I => \N__48752\
        );

    \I__11465\ : Span4Mux_s3_h
    port map (
            O => \N__48758\,
            I => \N__48749\
        );

    \I__11464\ : Span4Mux_s2_h
    port map (
            O => \N__48755\,
            I => \N__48746\
        );

    \I__11463\ : Sp12to4
    port map (
            O => \N__48752\,
            I => \N__48743\
        );

    \I__11462\ : Span4Mux_h
    port map (
            O => \N__48749\,
            I => \N__48740\
        );

    \I__11461\ : Span4Mux_h
    port map (
            O => \N__48746\,
            I => \N__48737\
        );

    \I__11460\ : Span12Mux_s11_h
    port map (
            O => \N__48743\,
            I => \N__48734\
        );

    \I__11459\ : Span4Mux_v
    port map (
            O => \N__48740\,
            I => \N__48731\
        );

    \I__11458\ : Span4Mux_h
    port map (
            O => \N__48737\,
            I => \N__48728\
        );

    \I__11457\ : Odrv12
    port map (
            O => \N__48734\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11456\ : Odrv4
    port map (
            O => \N__48731\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11455\ : Odrv4
    port map (
            O => \N__48728\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48717\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48713\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__48717\,
            I => \N__48710\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48716\,
            I => \N__48707\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__48713\,
            I => \N__48704\
        );

    \I__11449\ : Span4Mux_v
    port map (
            O => \N__48710\,
            I => \N__48701\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__48707\,
            I => \N__48698\
        );

    \I__11447\ : Odrv4
    port map (
            O => \N__48704\,
            I => pwm_duty_input_3
        );

    \I__11446\ : Odrv4
    port map (
            O => \N__48701\,
            I => pwm_duty_input_3
        );

    \I__11445\ : Odrv4
    port map (
            O => \N__48698\,
            I => pwm_duty_input_3
        );

    \I__11444\ : CascadeMux
    port map (
            O => \N__48691\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48688\,
            I => \N__48685\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__48685\,
            I => \N__48680\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48684\,
            I => \N__48675\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48675\
        );

    \I__11439\ : Odrv4
    port map (
            O => \N__48680\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__48675\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__11437\ : CascadeMux
    port map (
            O => \N__48670\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__11436\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48664\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48664\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48661\,
            I => \N__48658\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__48658\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__11432\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48652\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__48652\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48649\,
            I => \N__48644\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48648\,
            I => \N__48641\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48647\,
            I => \N__48638\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__48644\,
            I => \N__48635\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48641\,
            I => \N__48632\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48638\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__11424\ : Odrv12
    port map (
            O => \N__48635\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__11423\ : Odrv4
    port map (
            O => \N__48632\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48620\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48617\
        );

    \I__11420\ : CascadeMux
    port map (
            O => \N__48623\,
            I => \N__48614\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48620\,
            I => \N__48608\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48617\,
            I => \N__48608\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48614\,
            I => \N__48605\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48613\,
            I => \N__48602\
        );

    \I__11415\ : Span4Mux_v
    port map (
            O => \N__48608\,
            I => \N__48599\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48605\,
            I => \N__48596\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__48602\,
            I => \N__48593\
        );

    \I__11412\ : Span4Mux_h
    port map (
            O => \N__48599\,
            I => \N__48590\
        );

    \I__11411\ : Span4Mux_v
    port map (
            O => \N__48596\,
            I => \N__48587\
        );

    \I__11410\ : Odrv4
    port map (
            O => \N__48593\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__11409\ : Odrv4
    port map (
            O => \N__48590\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__11408\ : Odrv4
    port map (
            O => \N__48587\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48580\,
            I => \N__48574\
        );

    \I__11406\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48574\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48574\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__11404\ : CascadeMux
    port map (
            O => \N__48571\,
            I => \N__48567\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48564\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48561\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48564\,
            I => \N__48558\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48561\,
            I => \N__48555\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__48558\,
            I => \N__48551\
        );

    \I__11398\ : Span4Mux_h
    port map (
            O => \N__48555\,
            I => \N__48548\
        );

    \I__11397\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48545\
        );

    \I__11396\ : Span4Mux_h
    port map (
            O => \N__48551\,
            I => \N__48542\
        );

    \I__11395\ : Span4Mux_h
    port map (
            O => \N__48548\,
            I => \N__48539\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__48545\,
            I => \N__48536\
        );

    \I__11393\ : Span4Mux_h
    port map (
            O => \N__48542\,
            I => \N__48533\
        );

    \I__11392\ : Span4Mux_h
    port map (
            O => \N__48539\,
            I => \N__48530\
        );

    \I__11391\ : Span12Mux_h
    port map (
            O => \N__48536\,
            I => \N__48527\
        );

    \I__11390\ : Span4Mux_v
    port map (
            O => \N__48533\,
            I => \N__48522\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__48530\,
            I => \N__48522\
        );

    \I__11388\ : Odrv12
    port map (
            O => \N__48527\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__48522\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48517\,
            I => \N__48513\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48516\,
            I => \N__48510\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__48513\,
            I => \N__48507\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48504\
        );

    \I__11382\ : Span4Mux_h
    port map (
            O => \N__48507\,
            I => \N__48501\
        );

    \I__11381\ : Span4Mux_h
    port map (
            O => \N__48504\,
            I => \N__48498\
        );

    \I__11380\ : Span4Mux_h
    port map (
            O => \N__48501\,
            I => \N__48495\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__48498\,
            I => \N__48490\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__48495\,
            I => \N__48487\
        );

    \I__11377\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48482\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48482\
        );

    \I__11375\ : Span4Mux_h
    port map (
            O => \N__48490\,
            I => \N__48479\
        );

    \I__11374\ : Span4Mux_v
    port map (
            O => \N__48487\,
            I => \N__48476\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48482\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__11372\ : Odrv4
    port map (
            O => \N__48479\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__48476\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__11370\ : ClkMux
    port map (
            O => \N__48469\,
            I => \N__48466\
        );

    \I__11369\ : GlobalMux
    port map (
            O => \N__48466\,
            I => \N__48463\
        );

    \I__11368\ : gio2CtrlBuf
    port map (
            O => \N__48463\,
            I => delay_tr_input_c_g
        );

    \I__11367\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48455\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48459\,
            I => \N__48452\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48458\,
            I => \N__48449\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__48455\,
            I => \N__48446\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__48452\,
            I => \N__48443\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__48449\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__11361\ : Odrv12
    port map (
            O => \N__48446\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__11360\ : Odrv12
    port map (
            O => \N__48443\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__11359\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48433\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__48433\,
            I => \N__48428\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48425\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48422\
        );

    \I__11355\ : Span4Mux_v
    port map (
            O => \N__48428\,
            I => \N__48414\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48425\,
            I => \N__48414\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48414\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48411\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__48414\,
            I => \N__48406\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__48411\,
            I => \N__48406\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__48406\,
            I => \N__48403\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__48403\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__48400\,
            I => \N__48386\
        );

    \I__11346\ : InMux
    port map (
            O => \N__48399\,
            I => \N__48375\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48398\,
            I => \N__48375\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48397\,
            I => \N__48375\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48366\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48366\
        );

    \I__11341\ : InMux
    port map (
            O => \N__48394\,
            I => \N__48366\
        );

    \I__11340\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48366\
        );

    \I__11339\ : CascadeMux
    port map (
            O => \N__48392\,
            I => \N__48363\
        );

    \I__11338\ : CascadeMux
    port map (
            O => \N__48391\,
            I => \N__48359\
        );

    \I__11337\ : InMux
    port map (
            O => \N__48390\,
            I => \N__48339\
        );

    \I__11336\ : InMux
    port map (
            O => \N__48389\,
            I => \N__48339\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48386\,
            I => \N__48339\
        );

    \I__11334\ : InMux
    port map (
            O => \N__48385\,
            I => \N__48339\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48332\
        );

    \I__11332\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48332\
        );

    \I__11331\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48332\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48310\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48366\,
            I => \N__48310\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48303\
        );

    \I__11327\ : InMux
    port map (
            O => \N__48362\,
            I => \N__48303\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48359\,
            I => \N__48303\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48358\,
            I => \N__48300\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48357\,
            I => \N__48288\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48356\,
            I => \N__48288\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48355\,
            I => \N__48288\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48288\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48285\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48279\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48260\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48350\,
            I => \N__48260\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48260\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48257\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48339\,
            I => \N__48252\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__48332\,
            I => \N__48252\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48331\,
            I => \N__48247\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48247\
        );

    \I__11310\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48244\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48328\,
            I => \N__48239\
        );

    \I__11308\ : InMux
    port map (
            O => \N__48327\,
            I => \N__48224\
        );

    \I__11307\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48224\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48224\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48224\
        );

    \I__11304\ : InMux
    port map (
            O => \N__48323\,
            I => \N__48224\
        );

    \I__11303\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48224\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48321\,
            I => \N__48224\
        );

    \I__11301\ : InMux
    port map (
            O => \N__48320\,
            I => \N__48218\
        );

    \I__11300\ : InMux
    port map (
            O => \N__48319\,
            I => \N__48215\
        );

    \I__11299\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48210\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48317\,
            I => \N__48210\
        );

    \I__11297\ : InMux
    port map (
            O => \N__48316\,
            I => \N__48207\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48204\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__48310\,
            I => \N__48197\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__48303\,
            I => \N__48197\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__48300\,
            I => \N__48197\
        );

    \I__11292\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48194\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48191\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48297\,
            I => \N__48188\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__48288\,
            I => \N__48183\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__48285\,
            I => \N__48183\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48176\
        );

    \I__11286\ : InMux
    port map (
            O => \N__48283\,
            I => \N__48176\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48282\,
            I => \N__48176\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__48279\,
            I => \N__48149\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48144\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48144\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48141\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48138\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48135\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48126\
        );

    \I__11277\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48126\
        );

    \I__11276\ : InMux
    port map (
            O => \N__48271\,
            I => \N__48126\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48270\,
            I => \N__48126\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48269\,
            I => \N__48119\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48119\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48119\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__48260\,
            I => \N__48114\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__48257\,
            I => \N__48114\
        );

    \I__11269\ : Span4Mux_h
    port map (
            O => \N__48252\,
            I => \N__48111\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48106\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__48244\,
            I => \N__48106\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48101\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48101\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__48239\,
            I => \N__48096\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__48224\,
            I => \N__48096\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48223\,
            I => \N__48089\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48222\,
            I => \N__48089\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48221\,
            I => \N__48089\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48218\,
            I => \N__48084\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__48215\,
            I => \N__48084\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__48210\,
            I => \N__48081\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48207\,
            I => \N__48078\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__48204\,
            I => \N__48075\
        );

    \I__11254\ : Span4Mux_v
    port map (
            O => \N__48197\,
            I => \N__48072\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__48194\,
            I => \N__48061\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__48191\,
            I => \N__48061\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__48188\,
            I => \N__48061\
        );

    \I__11250\ : Span4Mux_v
    port map (
            O => \N__48183\,
            I => \N__48061\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48176\,
            I => \N__48061\
        );

    \I__11248\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48056\
        );

    \I__11247\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48056\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48049\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48172\,
            I => \N__48049\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48049\
        );

    \I__11243\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48044\
        );

    \I__11242\ : InMux
    port map (
            O => \N__48169\,
            I => \N__48044\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48035\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48167\,
            I => \N__48035\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48035\
        );

    \I__11238\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48035\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48164\,
            I => \N__48032\
        );

    \I__11236\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48017\
        );

    \I__11235\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48017\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48017\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48017\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48017\
        );

    \I__11231\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48017\
        );

    \I__11230\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48017\
        );

    \I__11229\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48014\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48007\
        );

    \I__11227\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48007\
        );

    \I__11226\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48007\
        );

    \I__11225\ : InMux
    port map (
            O => \N__48152\,
            I => \N__48004\
        );

    \I__11224\ : Span4Mux_h
    port map (
            O => \N__48149\,
            I => \N__47999\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__48144\,
            I => \N__47999\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__47996\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__48138\,
            I => \N__47985\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48135\,
            I => \N__47985\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__48126\,
            I => \N__47985\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__48119\,
            I => \N__47985\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__48114\,
            I => \N__47985\
        );

    \I__11216\ : Span4Mux_v
    port map (
            O => \N__48111\,
            I => \N__47980\
        );

    \I__11215\ : Span4Mux_h
    port map (
            O => \N__48106\,
            I => \N__47980\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__47961\
        );

    \I__11213\ : Span4Mux_v
    port map (
            O => \N__48096\,
            I => \N__47961\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__48089\,
            I => \N__47961\
        );

    \I__11211\ : Span4Mux_v
    port map (
            O => \N__48084\,
            I => \N__47961\
        );

    \I__11210\ : Span4Mux_v
    port map (
            O => \N__48081\,
            I => \N__47961\
        );

    \I__11209\ : Span4Mux_h
    port map (
            O => \N__48078\,
            I => \N__47961\
        );

    \I__11208\ : Span4Mux_v
    port map (
            O => \N__48075\,
            I => \N__47961\
        );

    \I__11207\ : Span4Mux_h
    port map (
            O => \N__48072\,
            I => \N__47961\
        );

    \I__11206\ : Span4Mux_v
    port map (
            O => \N__48061\,
            I => \N__47961\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48056\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__48049\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__48044\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__48035\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__48032\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__48017\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__48014\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__48007\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__48004\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11196\ : Odrv4
    port map (
            O => \N__47999\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11195\ : Odrv4
    port map (
            O => \N__47996\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11194\ : Odrv4
    port map (
            O => \N__47985\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11193\ : Odrv4
    port map (
            O => \N__47980\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11192\ : Odrv4
    port map (
            O => \N__47961\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11191\ : InMux
    port map (
            O => \N__47932\,
            I => \N__47928\
        );

    \I__11190\ : InMux
    port map (
            O => \N__47931\,
            I => \N__47925\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__47928\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__47925\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__11187\ : CEMux
    port map (
            O => \N__47920\,
            I => \N__47890\
        );

    \I__11186\ : CEMux
    port map (
            O => \N__47919\,
            I => \N__47890\
        );

    \I__11185\ : CEMux
    port map (
            O => \N__47918\,
            I => \N__47890\
        );

    \I__11184\ : CEMux
    port map (
            O => \N__47917\,
            I => \N__47890\
        );

    \I__11183\ : CEMux
    port map (
            O => \N__47916\,
            I => \N__47890\
        );

    \I__11182\ : CEMux
    port map (
            O => \N__47915\,
            I => \N__47890\
        );

    \I__11181\ : CEMux
    port map (
            O => \N__47914\,
            I => \N__47890\
        );

    \I__11180\ : CEMux
    port map (
            O => \N__47913\,
            I => \N__47890\
        );

    \I__11179\ : CEMux
    port map (
            O => \N__47912\,
            I => \N__47890\
        );

    \I__11178\ : CEMux
    port map (
            O => \N__47911\,
            I => \N__47890\
        );

    \I__11177\ : GlobalMux
    port map (
            O => \N__47890\,
            I => \N__47887\
        );

    \I__11176\ : gio2CtrlBuf
    port map (
            O => \N__47887\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__11175\ : InMux
    port map (
            O => \N__47884\,
            I => \N__47881\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__47881\,
            I => \N__47877\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47880\,
            I => \N__47874\
        );

    \I__11172\ : Span12Mux_v
    port map (
            O => \N__47877\,
            I => \N__47871\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__47874\,
            I => \N__47868\
        );

    \I__11170\ : Span12Mux_h
    port map (
            O => \N__47871\,
            I => \N__47863\
        );

    \I__11169\ : Span12Mux_s9_h
    port map (
            O => \N__47868\,
            I => \N__47863\
        );

    \I__11168\ : Odrv12
    port map (
            O => \N__47863\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47860\,
            I => \N__47857\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__47857\,
            I => \N__47854\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__47854\,
            I => \N__47851\
        );

    \I__11164\ : Odrv4
    port map (
            O => \N__47851\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__11163\ : InMux
    port map (
            O => \N__47848\,
            I => \N__47845\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__47845\,
            I => \N__47835\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47844\,
            I => \N__47820\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47820\
        );

    \I__11159\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47820\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47820\
        );

    \I__11157\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47820\
        );

    \I__11156\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47820\
        );

    \I__11155\ : InMux
    port map (
            O => \N__47838\,
            I => \N__47820\
        );

    \I__11154\ : Span4Mux_v
    port map (
            O => \N__47835\,
            I => \N__47813\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__47820\,
            I => \N__47813\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47819\,
            I => \N__47808\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47818\,
            I => \N__47808\
        );

    \I__11150\ : Span4Mux_v
    port map (
            O => \N__47813\,
            I => \N__47803\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47808\,
            I => \N__47803\
        );

    \I__11148\ : Span4Mux_h
    port map (
            O => \N__47803\,
            I => \N__47800\
        );

    \I__11147\ : Span4Mux_h
    port map (
            O => \N__47800\,
            I => \N__47797\
        );

    \I__11146\ : Odrv4
    port map (
            O => \N__47797\,
            I => \pwm_generator_inst.N_16\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__47794\,
            I => \N__47791\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47788\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47785\
        );

    \I__11142\ : Span4Mux_h
    port map (
            O => \N__47785\,
            I => \N__47782\
        );

    \I__11141\ : Odrv4
    port map (
            O => \N__47782\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__11140\ : CascadeMux
    port map (
            O => \N__47779\,
            I => \N__47776\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47776\,
            I => \N__47770\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47770\
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__47770\,
            I => \N__47766\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47769\,
            I => \N__47763\
        );

    \I__11135\ : Span4Mux_h
    port map (
            O => \N__47766\,
            I => \N__47760\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__47763\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__11133\ : Odrv4
    port map (
            O => \N__47760\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__11132\ : CascadeMux
    port map (
            O => \N__47755\,
            I => \N__47750\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47754\,
            I => \N__47747\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47742\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47750\,
            I => \N__47742\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__47747\,
            I => \N__47737\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47742\,
            I => \N__47737\
        );

    \I__11126\ : Odrv4
    port map (
            O => \N__47737\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47734\,
            I => \N__47731\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__47731\,
            I => \N__47728\
        );

    \I__11123\ : Span4Mux_h
    port map (
            O => \N__47728\,
            I => \N__47725\
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__47725\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__11121\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47719\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47719\,
            I => \N__47716\
        );

    \I__11119\ : Span4Mux_h
    port map (
            O => \N__47716\,
            I => \N__47712\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47715\,
            I => \N__47708\
        );

    \I__11117\ : Span4Mux_h
    port map (
            O => \N__47712\,
            I => \N__47705\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47702\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__47708\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__47705\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__47702\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47695\,
            I => \N__47690\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47694\,
            I => \N__47686\
        );

    \I__11110\ : CascadeMux
    port map (
            O => \N__47693\,
            I => \N__47683\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__47690\,
            I => \N__47680\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47677\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47686\,
            I => \N__47674\
        );

    \I__11106\ : InMux
    port map (
            O => \N__47683\,
            I => \N__47671\
        );

    \I__11105\ : Span4Mux_v
    port map (
            O => \N__47680\,
            I => \N__47668\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47677\,
            I => \N__47665\
        );

    \I__11103\ : Span4Mux_h
    port map (
            O => \N__47674\,
            I => \N__47662\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__47671\,
            I => \N__47659\
        );

    \I__11101\ : Span4Mux_h
    port map (
            O => \N__47668\,
            I => \N__47656\
        );

    \I__11100\ : Span4Mux_v
    port map (
            O => \N__47665\,
            I => \N__47651\
        );

    \I__11099\ : Span4Mux_h
    port map (
            O => \N__47662\,
            I => \N__47651\
        );

    \I__11098\ : Span4Mux_h
    port map (
            O => \N__47659\,
            I => \N__47648\
        );

    \I__11097\ : Odrv4
    port map (
            O => \N__47656\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__11096\ : Odrv4
    port map (
            O => \N__47651\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__47648\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47635\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47635\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47635\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47629\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47629\,
            I => \N__47626\
        );

    \I__11089\ : Span4Mux_h
    port map (
            O => \N__47626\,
            I => \N__47621\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47618\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47615\
        );

    \I__11086\ : Span4Mux_h
    port map (
            O => \N__47621\,
            I => \N__47612\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47609\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47615\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__47612\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__47609\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47602\,
            I => \N__47598\
        );

    \I__11080\ : InMux
    port map (
            O => \N__47601\,
            I => \N__47595\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47598\,
            I => \N__47590\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__47595\,
            I => \N__47587\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47584\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47581\
        );

    \I__11075\ : Span4Mux_h
    port map (
            O => \N__47590\,
            I => \N__47578\
        );

    \I__11074\ : Span4Mux_h
    port map (
            O => \N__47587\,
            I => \N__47575\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__47584\,
            I => \N__47572\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47581\,
            I => \N__47569\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__47578\,
            I => \N__47566\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__47575\,
            I => \N__47561\
        );

    \I__11069\ : Span4Mux_v
    port map (
            O => \N__47572\,
            I => \N__47561\
        );

    \I__11068\ : Odrv12
    port map (
            O => \N__47569\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11067\ : Odrv4
    port map (
            O => \N__47566\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__47561\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47548\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47553\,
            I => \N__47548\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__47548\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47545\,
            I => \N__47540\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47544\,
            I => \N__47537\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47534\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__47540\,
            I => \N__47531\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__47537\,
            I => \N__47528\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47534\,
            I => \N__47525\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__47531\,
            I => \N__47519\
        );

    \I__11055\ : Span4Mux_v
    port map (
            O => \N__47528\,
            I => \N__47519\
        );

    \I__11054\ : Span4Mux_v
    port map (
            O => \N__47525\,
            I => \N__47516\
        );

    \I__11053\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47513\
        );

    \I__11052\ : Span4Mux_h
    port map (
            O => \N__47519\,
            I => \N__47510\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__47516\,
            I => \N__47507\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47513\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__11049\ : Odrv4
    port map (
            O => \N__47510\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__11048\ : Odrv4
    port map (
            O => \N__47507\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__11047\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47497\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__47497\,
            I => \N__47493\
        );

    \I__11045\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47489\
        );

    \I__11044\ : Span4Mux_h
    port map (
            O => \N__47493\,
            I => \N__47486\
        );

    \I__11043\ : InMux
    port map (
            O => \N__47492\,
            I => \N__47483\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__47489\,
            I => \N__47480\
        );

    \I__11041\ : Span4Mux_h
    port map (
            O => \N__47486\,
            I => \N__47477\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47483\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__11039\ : Odrv4
    port map (
            O => \N__47480\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__11038\ : Odrv4
    port map (
            O => \N__47477\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__11037\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47467\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47467\,
            I => \N__47464\
        );

    \I__11035\ : Odrv4
    port map (
            O => \N__47464\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47455\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47455\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__47455\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__11031\ : CascadeMux
    port map (
            O => \N__47452\,
            I => \N__47448\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47442\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47448\,
            I => \N__47442\
        );

    \I__11028\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47439\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47436\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__47439\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__11025\ : Odrv4
    port map (
            O => \N__47436\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__11024\ : CascadeMux
    port map (
            O => \N__47431\,
            I => \N__47427\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47430\,
            I => \N__47421\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47427\,
            I => \N__47421\
        );

    \I__11021\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47418\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__47421\,
            I => \N__47415\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__47418\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__47415\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11017\ : CascadeMux
    port map (
            O => \N__47410\,
            I => \N__47407\
        );

    \I__11016\ : InMux
    port map (
            O => \N__47407\,
            I => \N__47404\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47401\
        );

    \I__11014\ : Odrv4
    port map (
            O => \N__47401\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47398\,
            I => \N__47394\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47397\,
            I => \N__47391\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__47394\,
            I => \N__47388\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__47391\,
            I => \N__47381\
        );

    \I__11009\ : Span4Mux_v
    port map (
            O => \N__47388\,
            I => \N__47381\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47387\,
            I => \N__47378\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47386\,
            I => \N__47375\
        );

    \I__11006\ : Span4Mux_h
    port map (
            O => \N__47381\,
            I => \N__47372\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__47378\,
            I => \N__47367\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__47375\,
            I => \N__47367\
        );

    \I__11003\ : Odrv4
    port map (
            O => \N__47372\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11002\ : Odrv4
    port map (
            O => \N__47367\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11001\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47359\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47359\,
            I => \N__47354\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47351\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47348\
        );

    \I__10997\ : Span4Mux_h
    port map (
            O => \N__47354\,
            I => \N__47345\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47351\,
            I => \N__47342\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__47348\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__10994\ : Odrv4
    port map (
            O => \N__47345\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__10993\ : Odrv12
    port map (
            O => \N__47342\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47335\,
            I => \N__47330\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47327\
        );

    \I__10990\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47324\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47330\,
            I => \N__47318\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47318\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__47324\,
            I => \N__47315\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47312\
        );

    \I__10985\ : Span4Mux_h
    port map (
            O => \N__47318\,
            I => \N__47309\
        );

    \I__10984\ : Span12Mux_s8_v
    port map (
            O => \N__47315\,
            I => \N__47306\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47312\,
            I => \N__47303\
        );

    \I__10982\ : Odrv4
    port map (
            O => \N__47309\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10981\ : Odrv12
    port map (
            O => \N__47306\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10980\ : Odrv4
    port map (
            O => \N__47303\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10979\ : InMux
    port map (
            O => \N__47296\,
            I => \N__47293\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47293\,
            I => \N__47288\
        );

    \I__10977\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47285\
        );

    \I__10976\ : InMux
    port map (
            O => \N__47291\,
            I => \N__47282\
        );

    \I__10975\ : Span4Mux_h
    port map (
            O => \N__47288\,
            I => \N__47277\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47285\,
            I => \N__47277\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__47282\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__10972\ : Odrv4
    port map (
            O => \N__47277\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__10971\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47267\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47264\
        );

    \I__10969\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47261\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__47267\,
            I => \N__47258\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47261\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__10965\ : Odrv4
    port map (
            O => \N__47258\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__10964\ : Odrv4
    port map (
            O => \N__47255\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47248\,
            I => \N__47245\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47245\,
            I => \N__47240\
        );

    \I__10961\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47237\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47234\
        );

    \I__10959\ : Span4Mux_v
    port map (
            O => \N__47240\,
            I => \N__47231\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47228\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__47234\,
            I => \N__47225\
        );

    \I__10956\ : Span4Mux_h
    port map (
            O => \N__47231\,
            I => \N__47221\
        );

    \I__10955\ : Span4Mux_v
    port map (
            O => \N__47228\,
            I => \N__47216\
        );

    \I__10954\ : Span4Mux_v
    port map (
            O => \N__47225\,
            I => \N__47216\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47213\
        );

    \I__10952\ : Odrv4
    port map (
            O => \N__47221\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__10951\ : Odrv4
    port map (
            O => \N__47216\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__47213\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__10949\ : InMux
    port map (
            O => \N__47206\,
            I => \N__47203\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47203\,
            I => \N__47200\
        );

    \I__10947\ : Span4Mux_h
    port map (
            O => \N__47200\,
            I => \N__47197\
        );

    \I__10946\ : Odrv4
    port map (
            O => \N__47197\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47191\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47186\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47181\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47181\
        );

    \I__10941\ : Span4Mux_v
    port map (
            O => \N__47186\,
            I => \N__47177\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47181\,
            I => \N__47174\
        );

    \I__10939\ : CascadeMux
    port map (
            O => \N__47180\,
            I => \N__47171\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__47177\,
            I => \N__47166\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__47174\,
            I => \N__47166\
        );

    \I__10936\ : InMux
    port map (
            O => \N__47171\,
            I => \N__47163\
        );

    \I__10935\ : Odrv4
    port map (
            O => \N__47166\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47163\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10933\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47155\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47155\,
            I => \N__47151\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47148\
        );

    \I__10930\ : Odrv12
    port map (
            O => \N__47151\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47148\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47143\,
            I => \N__47140\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47140\,
            I => \N__47137\
        );

    \I__10926\ : Span4Mux_h
    port map (
            O => \N__47137\,
            I => \N__47134\
        );

    \I__10925\ : Odrv4
    port map (
            O => \N__47134\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__10924\ : CascadeMux
    port map (
            O => \N__47131\,
            I => \N__47128\
        );

    \I__10923\ : InMux
    port map (
            O => \N__47128\,
            I => \N__47123\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47120\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47117\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__47123\,
            I => \N__47112\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47112\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__47117\,
            I => \N__47107\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__47112\,
            I => \N__47107\
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__47107\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47104\,
            I => \N__47100\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47097\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47094\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47097\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__10911\ : Odrv4
    port map (
            O => \N__47094\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__47089\,
            I => \N__47085\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47082\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47085\,
            I => \N__47079\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__47082\,
            I => \N__47075\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__47079\,
            I => \N__47072\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47069\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__47075\,
            I => \N__47064\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__47072\,
            I => \N__47064\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__47069\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__47064\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10900\ : CascadeMux
    port map (
            O => \N__47059\,
            I => \N__47056\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47053\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47050\
        );

    \I__10897\ : Span4Mux_h
    port map (
            O => \N__47050\,
            I => \N__47047\
        );

    \I__10896\ : Span4Mux_h
    port map (
            O => \N__47047\,
            I => \N__47044\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__47044\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47041\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47038\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__10892\ : InMux
    port map (
            O => \N__47035\,
            I => \N__47031\
        );

    \I__10891\ : InMux
    port map (
            O => \N__47034\,
            I => \N__47027\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__47031\,
            I => \N__47024\
        );

    \I__10889\ : InMux
    port map (
            O => \N__47030\,
            I => \N__47021\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__47027\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__47024\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__47021\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47014\,
            I => \N__47011\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__47011\,
            I => \N__47007\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47010\,
            I => \N__47004\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__47007\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__47004\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10880\ : CascadeMux
    port map (
            O => \N__46999\,
            I => \N__46996\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46993\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__46993\,
            I => \N__46990\
        );

    \I__10877\ : Odrv12
    port map (
            O => \N__46990\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46983\
        );

    \I__10875\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46980\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46983\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__46980\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46972\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46972\,
            I => \N__46969\
        );

    \I__10870\ : Span4Mux_h
    port map (
            O => \N__46969\,
            I => \N__46962\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46959\
        );

    \I__10868\ : InMux
    port map (
            O => \N__46967\,
            I => \N__46956\
        );

    \I__10867\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46951\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46951\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__46962\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46959\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46956\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__46951\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46936\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46941\,
            I => \N__46931\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46931\
        );

    \I__10858\ : CascadeMux
    port map (
            O => \N__46939\,
            I => \N__46928\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__46936\,
            I => \N__46923\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46931\,
            I => \N__46923\
        );

    \I__10855\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46920\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__46923\,
            I => \N__46917\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__46920\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__10852\ : Odrv4
    port map (
            O => \N__46917\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__10851\ : CascadeMux
    port map (
            O => \N__46912\,
            I => \N__46908\
        );

    \I__10850\ : CascadeMux
    port map (
            O => \N__46911\,
            I => \N__46905\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46899\
        );

    \I__10848\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46896\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46904\,
            I => \N__46891\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46891\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46902\,
            I => \N__46888\
        );

    \I__10844\ : LocalMux
    port map (
            O => \N__46899\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46896\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__46891\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46888\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__10840\ : IoInMux
    port map (
            O => \N__46879\,
            I => \N__46876\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46876\,
            I => \N__46873\
        );

    \I__10838\ : IoSpan4Mux
    port map (
            O => \N__46873\,
            I => \N__46862\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46853\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46853\
        );

    \I__10835\ : InMux
    port map (
            O => \N__46870\,
            I => \N__46853\
        );

    \I__10834\ : InMux
    port map (
            O => \N__46869\,
            I => \N__46853\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46868\,
            I => \N__46846\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46846\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46846\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46865\,
            I => \N__46839\
        );

    \I__10829\ : Span4Mux_s3_v
    port map (
            O => \N__46862\,
            I => \N__46817\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46853\,
            I => \N__46812\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46812\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46845\,
            I => \N__46803\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46844\,
            I => \N__46803\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46843\,
            I => \N__46803\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46842\,
            I => \N__46803\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46839\,
            I => \N__46800\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46838\,
            I => \N__46793\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46793\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46836\,
            I => \N__46793\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46784\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46784\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46784\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46784\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46775\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46830\,
            I => \N__46775\
        );

    \I__10812\ : InMux
    port map (
            O => \N__46829\,
            I => \N__46775\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46775\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46766\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46826\,
            I => \N__46766\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46766\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46766\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46757\
        );

    \I__10805\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46757\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46757\
        );

    \I__10803\ : InMux
    port map (
            O => \N__46820\,
            I => \N__46757\
        );

    \I__10802\ : Sp12to4
    port map (
            O => \N__46817\,
            I => \N__46754\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__46812\,
            I => \N__46747\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__46803\,
            I => \N__46747\
        );

    \I__10799\ : Span4Mux_h
    port map (
            O => \N__46800\,
            I => \N__46747\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46793\,
            I => \N__46736\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__46784\,
            I => \N__46736\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__46775\,
            I => \N__46736\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__46766\,
            I => \N__46736\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__46757\,
            I => \N__46736\
        );

    \I__10793\ : Span12Mux_v
    port map (
            O => \N__46754\,
            I => \N__46733\
        );

    \I__10792\ : Odrv4
    port map (
            O => \N__46747\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10791\ : Odrv12
    port map (
            O => \N__46736\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10790\ : Odrv12
    port map (
            O => \N__46733\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46726\,
            I => \N__46723\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46723\,
            I => \N__46719\
        );

    \I__10787\ : InMux
    port map (
            O => \N__46722\,
            I => \N__46716\
        );

    \I__10786\ : Span4Mux_h
    port map (
            O => \N__46719\,
            I => \N__46713\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__46716\,
            I => \N__46710\
        );

    \I__10784\ : Span4Mux_h
    port map (
            O => \N__46713\,
            I => \N__46707\
        );

    \I__10783\ : Span4Mux_s3_h
    port map (
            O => \N__46710\,
            I => \N__46704\
        );

    \I__10782\ : Span4Mux_h
    port map (
            O => \N__46707\,
            I => \N__46699\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__46704\,
            I => \N__46699\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__46699\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46692\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46689\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46692\,
            I => \N__46684\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46689\,
            I => \N__46684\
        );

    \I__10775\ : Span4Mux_v
    port map (
            O => \N__46684\,
            I => \N__46681\
        );

    \I__10774\ : Odrv4
    port map (
            O => \N__46681\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46675\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46671\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46674\,
            I => \N__46668\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__46671\,
            I => \N__46663\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__46668\,
            I => \N__46663\
        );

    \I__10768\ : Span4Mux_h
    port map (
            O => \N__46663\,
            I => \N__46660\
        );

    \I__10767\ : Span4Mux_h
    port map (
            O => \N__46660\,
            I => \N__46657\
        );

    \I__10766\ : Odrv4
    port map (
            O => \N__46657\,
            I => \pwm_generator_inst.O_10\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46650\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46653\,
            I => \N__46646\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46650\,
            I => \N__46643\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46640\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__46646\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10760\ : Odrv12
    port map (
            O => \N__46643\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46640\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10758\ : IoInMux
    port map (
            O => \N__46633\,
            I => \N__46630\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__46630\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46620\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46626\,
            I => \N__46620\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46625\,
            I => \N__46617\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__46620\,
            I => \N__46614\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46617\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__10751\ : Odrv4
    port map (
            O => \N__46614\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46609\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__10749\ : CascadeMux
    port map (
            O => \N__46606\,
            I => \N__46602\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46597\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46597\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__46597\,
            I => \N__46593\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46596\,
            I => \N__46590\
        );

    \I__10744\ : Span4Mux_h
    port map (
            O => \N__46593\,
            I => \N__46587\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46590\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__10742\ : Odrv4
    port map (
            O => \N__46587\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46582\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46579\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46576\,
            I => \bfn_18_13_0_\
        );

    \I__10738\ : CascadeMux
    port map (
            O => \N__46573\,
            I => \N__46570\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46563\
        );

    \I__10736\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46563\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46568\,
            I => \N__46560\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46563\,
            I => \N__46557\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46560\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10732\ : Odrv12
    port map (
            O => \N__46557\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46552\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46549\,
            I => \N__46542\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46548\,
            I => \N__46542\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46539\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46536\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__46539\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10725\ : Odrv4
    port map (
            O => \N__46536\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46531\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__10723\ : CascadeMux
    port map (
            O => \N__46528\,
            I => \N__46525\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46520\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46517\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46514\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__46520\,
            I => \N__46511\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46517\,
            I => \N__46508\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46514\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10716\ : Odrv12
    port map (
            O => \N__46511\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10715\ : Odrv4
    port map (
            O => \N__46508\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10714\ : InMux
    port map (
            O => \N__46501\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46493\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46497\,
            I => \N__46490\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46496\,
            I => \N__46487\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__46493\,
            I => \N__46482\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__46490\,
            I => \N__46482\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__46487\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__46482\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10706\ : InMux
    port map (
            O => \N__46477\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46470\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46467\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46470\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__46467\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46462\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46455\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46452\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__46455\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__46452\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46447\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__10695\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46440\
        );

    \I__10694\ : InMux
    port map (
            O => \N__46443\,
            I => \N__46437\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__46440\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__46437\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46432\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__10690\ : InMux
    port map (
            O => \N__46429\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46426\,
            I => \bfn_18_12_0_\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__46423\,
            I => \N__46420\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46420\,
            I => \N__46415\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46419\,
            I => \N__46412\
        );

    \I__10685\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46409\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__46415\,
            I => \N__46406\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__46412\,
            I => \N__46403\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46409\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__46406\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10680\ : Odrv12
    port map (
            O => \N__46403\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10679\ : InMux
    port map (
            O => \N__46396\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__10678\ : CascadeMux
    port map (
            O => \N__46393\,
            I => \N__46389\
        );

    \I__10677\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46385\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46382\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46379\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__46385\,
            I => \N__46376\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__46382\,
            I => \N__46373\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46379\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10671\ : Odrv4
    port map (
            O => \N__46376\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10670\ : Odrv12
    port map (
            O => \N__46373\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46366\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__10668\ : CascadeMux
    port map (
            O => \N__46363\,
            I => \N__46360\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46360\,
            I => \N__46355\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46352\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46349\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__46355\,
            I => \N__46344\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__46352\,
            I => \N__46344\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__46349\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__46344\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__10660\ : InMux
    port map (
            O => \N__46339\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46331\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46328\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46334\,
            I => \N__46325\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46331\,
            I => \N__46320\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46328\,
            I => \N__46320\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46325\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__46320\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46315\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__10651\ : InMux
    port map (
            O => \N__46312\,
            I => \N__46308\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46311\,
            I => \N__46305\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__46308\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__46305\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46300\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46293\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46290\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__46293\,
            I => \N__46287\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46290\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10642\ : Odrv4
    port map (
            O => \N__46287\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46282\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__10640\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46275\
        );

    \I__10639\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46272\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46275\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46272\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46267\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46260\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46263\,
            I => \N__46257\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46254\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46257\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10631\ : Odrv4
    port map (
            O => \N__46254\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10630\ : InMux
    port map (
            O => \N__46249\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__10629\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46242\
        );

    \I__10628\ : InMux
    port map (
            O => \N__46245\,
            I => \N__46239\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46242\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__46239\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10625\ : InMux
    port map (
            O => \N__46234\,
            I => \bfn_18_11_0_\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46227\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46230\,
            I => \N__46224\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__46227\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__46224\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46219\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46216\,
            I => \N__46212\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46215\,
            I => \N__46209\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__46212\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__46209\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46204\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46197\
        );

    \I__10613\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46194\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__46197\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46194\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10610\ : InMux
    port map (
            O => \N__46189\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46186\,
            I => \N__46182\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46185\,
            I => \N__46178\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__46182\,
            I => \N__46175\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46172\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46178\,
            I => \N__46169\
        );

    \I__10604\ : Span4Mux_v
    port map (
            O => \N__46175\,
            I => \N__46163\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__46172\,
            I => \N__46163\
        );

    \I__10602\ : Span4Mux_v
    port map (
            O => \N__46169\,
            I => \N__46160\
        );

    \I__10601\ : InMux
    port map (
            O => \N__46168\,
            I => \N__46157\
        );

    \I__10600\ : Span4Mux_h
    port map (
            O => \N__46163\,
            I => \N__46154\
        );

    \I__10599\ : Odrv4
    port map (
            O => \N__46160\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__46157\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__46154\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46143\
        );

    \I__10595\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46140\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46137\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__46133\
        );

    \I__10592\ : Span4Mux_h
    port map (
            O => \N__46137\,
            I => \N__46130\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46127\
        );

    \I__10590\ : Span4Mux_h
    port map (
            O => \N__46133\,
            I => \N__46124\
        );

    \I__10589\ : Span4Mux_v
    port map (
            O => \N__46130\,
            I => \N__46121\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__46127\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10587\ : Odrv4
    port map (
            O => \N__46124\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10586\ : Odrv4
    port map (
            O => \N__46121\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10585\ : InMux
    port map (
            O => \N__46114\,
            I => \N__46111\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46111\,
            I => \N__46107\
        );

    \I__10583\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46104\
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__46107\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46104\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__46099\,
            I => \N__46095\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46092\
        );

    \I__10578\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46089\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__46092\,
            I => \N__46086\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46089\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__10575\ : Odrv4
    port map (
            O => \N__46086\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__10574\ : CascadeMux
    port map (
            O => \N__46081\,
            I => \N__46078\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46075\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__10571\ : Span4Mux_v
    port map (
            O => \N__46072\,
            I => \N__46069\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__46069\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__10569\ : InMux
    port map (
            O => \N__46066\,
            I => \N__46062\
        );

    \I__10568\ : InMux
    port map (
            O => \N__46065\,
            I => \N__46059\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__46062\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__46059\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__10565\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46050\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46047\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__46050\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__46047\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46042\,
            I => \N__46039\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__46039\,
            I => \N__46036\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__46036\,
            I => \N__46033\
        );

    \I__10558\ : Odrv4
    port map (
            O => \N__46033\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__10557\ : CascadeMux
    port map (
            O => \N__46030\,
            I => \N__46026\
        );

    \I__10556\ : InMux
    port map (
            O => \N__46029\,
            I => \N__46023\
        );

    \I__10555\ : InMux
    port map (
            O => \N__46026\,
            I => \N__46020\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46023\,
            I => \N__46017\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__46020\,
            I => \N__46011\
        );

    \I__10552\ : Span4Mux_v
    port map (
            O => \N__46017\,
            I => \N__46011\
        );

    \I__10551\ : InMux
    port map (
            O => \N__46016\,
            I => \N__46008\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__46011\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__46008\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10548\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45999\
        );

    \I__10547\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45996\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45999\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__45996\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45991\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__10543\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45985\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45985\,
            I => \N__45982\
        );

    \I__10541\ : Span4Mux_h
    port map (
            O => \N__45982\,
            I => \N__45979\
        );

    \I__10540\ : Odrv4
    port map (
            O => \N__45979\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__45976\,
            I => \N__45973\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45973\,
            I => \N__45969\
        );

    \I__10537\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45966\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__45969\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__45966\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45961\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45954\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45951\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45954\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__45951\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45946\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__45943\,
            I => \N__45938\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45935\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45932\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45938\,
            I => \N__45929\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45935\,
            I => \N__45925\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__45932\,
            I => \N__45922\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__45929\,
            I => \N__45919\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45928\,
            I => \N__45916\
        );

    \I__10520\ : Span4Mux_h
    port map (
            O => \N__45925\,
            I => \N__45913\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__45922\,
            I => \N__45908\
        );

    \I__10518\ : Span4Mux_v
    port map (
            O => \N__45919\,
            I => \N__45908\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__45916\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10516\ : Odrv4
    port map (
            O => \N__45913\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__45908\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45901\,
            I => \N__45897\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45894\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45890\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45894\,
            I => \N__45887\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45884\
        );

    \I__10509\ : Span4Mux_v
    port map (
            O => \N__45890\,
            I => \N__45881\
        );

    \I__10508\ : Span4Mux_v
    port map (
            O => \N__45887\,
            I => \N__45878\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45884\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10506\ : Odrv4
    port map (
            O => \N__45881\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10505\ : Odrv4
    port map (
            O => \N__45878\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45865\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45865\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__45865\,
            I => \N__45862\
        );

    \I__10501\ : Odrv4
    port map (
            O => \N__45862\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__45859\,
            I => \N__45856\
        );

    \I__10499\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10498\ : InMux
    port map (
            O => \N__45855\,
            I => \N__45850\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45847\
        );

    \I__10496\ : Odrv4
    port map (
            O => \N__45847\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__10495\ : CEMux
    port map (
            O => \N__45844\,
            I => \N__45841\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45841\,
            I => \N__45837\
        );

    \I__10493\ : CEMux
    port map (
            O => \N__45840\,
            I => \N__45829\
        );

    \I__10492\ : Span4Mux_h
    port map (
            O => \N__45837\,
            I => \N__45820\
        );

    \I__10491\ : CEMux
    port map (
            O => \N__45836\,
            I => \N__45817\
        );

    \I__10490\ : CEMux
    port map (
            O => \N__45835\,
            I => \N__45811\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45804\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45804\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45832\,
            I => \N__45804\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45829\,
            I => \N__45801\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45828\,
            I => \N__45798\
        );

    \I__10484\ : CEMux
    port map (
            O => \N__45827\,
            I => \N__45794\
        );

    \I__10483\ : CEMux
    port map (
            O => \N__45826\,
            I => \N__45791\
        );

    \I__10482\ : CEMux
    port map (
            O => \N__45825\,
            I => \N__45788\
        );

    \I__10481\ : CEMux
    port map (
            O => \N__45824\,
            I => \N__45785\
        );

    \I__10480\ : CEMux
    port map (
            O => \N__45823\,
            I => \N__45766\
        );

    \I__10479\ : Span4Mux_v
    port map (
            O => \N__45820\,
            I => \N__45761\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45761\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45816\,
            I => \N__45746\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45815\,
            I => \N__45746\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45814\,
            I => \N__45746\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45743\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45804\,
            I => \N__45736\
        );

    \I__10472\ : Span4Mux_h
    port map (
            O => \N__45801\,
            I => \N__45736\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__45798\,
            I => \N__45736\
        );

    \I__10470\ : CEMux
    port map (
            O => \N__45797\,
            I => \N__45733\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__45794\,
            I => \N__45726\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45791\,
            I => \N__45726\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45788\,
            I => \N__45726\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45785\,
            I => \N__45723\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45714\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45714\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45714\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45714\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45780\,
            I => \N__45705\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45705\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45705\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45777\,
            I => \N__45705\
        );

    \I__10457\ : InMux
    port map (
            O => \N__45776\,
            I => \N__45696\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45775\,
            I => \N__45696\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45696\
        );

    \I__10454\ : InMux
    port map (
            O => \N__45773\,
            I => \N__45696\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45772\,
            I => \N__45687\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45771\,
            I => \N__45687\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45770\,
            I => \N__45687\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45769\,
            I => \N__45687\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45766\,
            I => \N__45682\
        );

    \I__10448\ : Span4Mux_h
    port map (
            O => \N__45761\,
            I => \N__45682\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45760\,
            I => \N__45673\
        );

    \I__10446\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45673\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45673\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45673\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45664\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45664\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45754\,
            I => \N__45664\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45753\,
            I => \N__45664\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45746\,
            I => \N__45657\
        );

    \I__10438\ : Span4Mux_v
    port map (
            O => \N__45743\,
            I => \N__45657\
        );

    \I__10437\ : Span4Mux_v
    port map (
            O => \N__45736\,
            I => \N__45657\
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__45733\,
            I => \N__45650\
        );

    \I__10435\ : Sp12to4
    port map (
            O => \N__45726\,
            I => \N__45650\
        );

    \I__10434\ : Sp12to4
    port map (
            O => \N__45723\,
            I => \N__45650\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45714\,
            I => \N__45639\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45639\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45639\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45687\,
            I => \N__45639\
        );

    \I__10429\ : Span4Mux_v
    port map (
            O => \N__45682\,
            I => \N__45639\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45673\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45664\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__45657\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10425\ : Odrv12
    port map (
            O => \N__45650\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__45639\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__45628\,
            I => \N__45625\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45622\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45619\
        );

    \I__10420\ : Sp12to4
    port map (
            O => \N__45619\,
            I => \N__45616\
        );

    \I__10419\ : Odrv12
    port map (
            O => \N__45616\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45610\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45607\
        );

    \I__10416\ : Span4Mux_h
    port map (
            O => \N__45607\,
            I => \N__45602\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45599\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45596\
        );

    \I__10413\ : Span4Mux_v
    port map (
            O => \N__45602\,
            I => \N__45593\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45590\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45596\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10410\ : Odrv4
    port map (
            O => \N__45593\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10409\ : Odrv4
    port map (
            O => \N__45590\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45579\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45582\,
            I => \N__45575\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__45579\,
            I => \N__45571\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45568\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45575\,
            I => \N__45565\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45562\
        );

    \I__10402\ : Span4Mux_v
    port map (
            O => \N__45571\,
            I => \N__45557\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45568\,
            I => \N__45557\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__45565\,
            I => \N__45554\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__45562\,
            I => \N__45551\
        );

    \I__10398\ : Span4Mux_h
    port map (
            O => \N__45557\,
            I => \N__45548\
        );

    \I__10397\ : Odrv4
    port map (
            O => \N__45554\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10396\ : Odrv12
    port map (
            O => \N__45551\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__45548\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10394\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45538\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__45538\,
            I => \N__45533\
        );

    \I__10392\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45530\
        );

    \I__10391\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45527\
        );

    \I__10390\ : Span4Mux_h
    port map (
            O => \N__45533\,
            I => \N__45524\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45530\,
            I => \N__45521\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45527\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10387\ : Odrv4
    port map (
            O => \N__45524\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10386\ : Odrv4
    port map (
            O => \N__45521\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45510\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45506\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__45510\,
            I => \N__45503\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45499\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__45506\,
            I => \N__45496\
        );

    \I__10380\ : Span4Mux_v
    port map (
            O => \N__45503\,
            I => \N__45493\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45490\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45499\,
            I => \N__45487\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__45496\,
            I => \N__45484\
        );

    \I__10376\ : Odrv4
    port map (
            O => \N__45493\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__45490\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45487\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__45484\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10372\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45472\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45468\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45464\
        );

    \I__10369\ : Span4Mux_v
    port map (
            O => \N__45468\,
            I => \N__45461\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45467\,
            I => \N__45458\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__45464\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__10366\ : Odrv4
    port map (
            O => \N__45461\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__45458\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45447\
        );

    \I__10363\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45443\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__45447\,
            I => \N__45439\
        );

    \I__10361\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45436\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__45443\,
            I => \N__45433\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45430\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__45439\,
            I => \N__45427\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__45436\,
            I => \N__45422\
        );

    \I__10356\ : Span4Mux_v
    port map (
            O => \N__45433\,
            I => \N__45422\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__45430\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__10354\ : Odrv4
    port map (
            O => \N__45427\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__10353\ : Odrv4
    port map (
            O => \N__45422\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__45415\,
            I => \N__45412\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45409\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45409\,
            I => \N__45406\
        );

    \I__10349\ : Odrv4
    port map (
            O => \N__45406\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__45400\,
            I => \N__45394\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45391\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45388\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45385\
        );

    \I__10343\ : Span4Mux_v
    port map (
            O => \N__45394\,
            I => \N__45378\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__45391\,
            I => \N__45378\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__45388\,
            I => \N__45378\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__45385\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10339\ : Odrv4
    port map (
            O => \N__45378\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45373\,
            I => \N__45370\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__45370\,
            I => \N__45366\
        );

    \I__10336\ : InMux
    port map (
            O => \N__45369\,
            I => \N__45362\
        );

    \I__10335\ : Span4Mux_v
    port map (
            O => \N__45366\,
            I => \N__45359\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45365\,
            I => \N__45356\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__45362\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10332\ : Odrv4
    port map (
            O => \N__45359\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45356\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45346\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__45346\,
            I => \N__45343\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__45343\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45337\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45333\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45329\
        );

    \I__10324\ : Span4Mux_v
    port map (
            O => \N__45333\,
            I => \N__45326\
        );

    \I__10323\ : InMux
    port map (
            O => \N__45332\,
            I => \N__45323\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45329\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__10321\ : Odrv4
    port map (
            O => \N__45326\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45323\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45313\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__45313\,
            I => \N__45310\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__45310\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__10316\ : InMux
    port map (
            O => \N__45307\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45304\,
            I => \N__45301\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__45301\,
            I => \N__45297\
        );

    \I__10313\ : InMux
    port map (
            O => \N__45300\,
            I => \N__45293\
        );

    \I__10312\ : Span4Mux_v
    port map (
            O => \N__45297\,
            I => \N__45290\
        );

    \I__10311\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45287\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__45293\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__45290\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__45287\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45277\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__45277\,
            I => \N__45274\
        );

    \I__10305\ : Odrv4
    port map (
            O => \N__45274\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45271\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45268\,
            I => \N__45264\
        );

    \I__10302\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45261\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__45264\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45261\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45256\,
            I => \N__45253\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__45253\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45250\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45244\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__45244\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45241\,
            I => \bfn_17_28_0_\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45235\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45231\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45228\
        );

    \I__10290\ : Span4Mux_s3_v
    port map (
            O => \N__45231\,
            I => \N__45225\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45228\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45225\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45217\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45217\,
            I => \N__45214\
        );

    \I__10285\ : Span4Mux_v
    port map (
            O => \N__45214\,
            I => \N__45211\
        );

    \I__10284\ : Span4Mux_s2_v
    port map (
            O => \N__45211\,
            I => \N__45208\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__45208\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45205\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45197\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45194\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45191\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__45188\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45194\,
            I => \N__45185\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__45191\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__10275\ : Odrv4
    port map (
            O => \N__45188\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__10274\ : Odrv4
    port map (
            O => \N__45185\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45178\,
            I => \N__45175\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__45175\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__10271\ : InMux
    port map (
            O => \N__45172\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45169\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__10269\ : InMux
    port map (
            O => \N__45166\,
            I => \N__45163\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__45163\,
            I => \N__45160\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__45160\,
            I => \N__45157\
        );

    \I__10266\ : Odrv4
    port map (
            O => \N__45157\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__10265\ : CascadeMux
    port map (
            O => \N__45154\,
            I => \N__45150\
        );

    \I__10264\ : InMux
    port map (
            O => \N__45153\,
            I => \N__45147\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45144\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__45147\,
            I => \N__45141\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__45144\,
            I => \N__45138\
        );

    \I__10260\ : Span4Mux_h
    port map (
            O => \N__45141\,
            I => \N__45135\
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__45138\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__10258\ : Odrv4
    port map (
            O => \N__45135\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45125\
        );

    \I__10256\ : InMux
    port map (
            O => \N__45129\,
            I => \N__45120\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45120\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__45125\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__45120\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45115\,
            I => \N__45112\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__45112\,
            I => \N__45109\
        );

    \I__10250\ : Span4Mux_h
    port map (
            O => \N__45109\,
            I => \N__45106\
        );

    \I__10249\ : Span4Mux_h
    port map (
            O => \N__45106\,
            I => \N__45103\
        );

    \I__10248\ : Odrv4
    port map (
            O => \N__45103\,
            I => \pwm_generator_inst.O_5\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45097\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__45097\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45094\,
            I => \N__45091\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__45091\,
            I => \N__45088\
        );

    \I__10243\ : Span4Mux_h
    port map (
            O => \N__45088\,
            I => \N__45085\
        );

    \I__10242\ : Span4Mux_h
    port map (
            O => \N__45085\,
            I => \N__45082\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__45082\,
            I => \pwm_generator_inst.O_6\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45076\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__45076\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45073\,
            I => \N__45070\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__45070\,
            I => \N__45067\
        );

    \I__10236\ : Span4Mux_h
    port map (
            O => \N__45067\,
            I => \N__45064\
        );

    \I__10235\ : Span4Mux_h
    port map (
            O => \N__45064\,
            I => \N__45061\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__45061\,
            I => \pwm_generator_inst.O_7\
        );

    \I__10233\ : InMux
    port map (
            O => \N__45058\,
            I => \N__45055\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__45055\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__10231\ : InMux
    port map (
            O => \N__45052\,
            I => \N__45049\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__45049\,
            I => \N__45046\
        );

    \I__10229\ : Span4Mux_v
    port map (
            O => \N__45046\,
            I => \N__45043\
        );

    \I__10228\ : Span4Mux_h
    port map (
            O => \N__45043\,
            I => \N__45040\
        );

    \I__10227\ : Span4Mux_h
    port map (
            O => \N__45040\,
            I => \N__45037\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__45037\,
            I => \pwm_generator_inst.O_8\
        );

    \I__10225\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45031\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__45031\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45028\,
            I => \N__45025\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__45025\,
            I => \N__45022\
        );

    \I__10221\ : Span4Mux_v
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__10220\ : Span4Mux_h
    port map (
            O => \N__45019\,
            I => \N__45016\
        );

    \I__10219\ : Span4Mux_h
    port map (
            O => \N__45016\,
            I => \N__45013\
        );

    \I__10218\ : Odrv4
    port map (
            O => \N__45013\,
            I => \pwm_generator_inst.O_9\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45007\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__45007\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__10215\ : InMux
    port map (
            O => \N__45004\,
            I => \N__45001\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44998\
        );

    \I__10213\ : Odrv12
    port map (
            O => \N__44998\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__10212\ : InMux
    port map (
            O => \N__44995\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__44992\,
            I => \N__44986\
        );

    \I__10210\ : CascadeMux
    port map (
            O => \N__44991\,
            I => \N__44980\
        );

    \I__10209\ : CascadeMux
    port map (
            O => \N__44990\,
            I => \N__44977\
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__44989\,
            I => \N__44973\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44968\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44961\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44961\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44961\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44956\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44956\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44953\
        );

    \I__10200\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44950\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__44972\,
            I => \N__44946\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44942\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44968\,
            I => \N__44937\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44937\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__44956\,
            I => \N__44934\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44929\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44929\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44926\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44921\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44921\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__44942\,
            I => \N__44918\
        );

    \I__10188\ : Span4Mux_h
    port map (
            O => \N__44937\,
            I => \N__44913\
        );

    \I__10187\ : Span4Mux_h
    port map (
            O => \N__44934\,
            I => \N__44913\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__44929\,
            I => \N__44908\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__44926\,
            I => \N__44908\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__44921\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__44918\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__44913\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__10181\ : Odrv4
    port map (
            O => \N__44908\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44895\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44892\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44889\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44886\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__44889\,
            I => \N__44883\
        );

    \I__10175\ : Span4Mux_h
    port map (
            O => \N__44886\,
            I => \N__44880\
        );

    \I__10174\ : Span4Mux_h
    port map (
            O => \N__44883\,
            I => \N__44877\
        );

    \I__10173\ : Span4Mux_h
    port map (
            O => \N__44880\,
            I => \N__44874\
        );

    \I__10172\ : Span4Mux_h
    port map (
            O => \N__44877\,
            I => \N__44871\
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__44874\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__10170\ : Odrv4
    port map (
            O => \N__44871\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44863\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44863\,
            I => \N__44860\
        );

    \I__10167\ : Span4Mux_h
    port map (
            O => \N__44860\,
            I => \N__44857\
        );

    \I__10166\ : Odrv4
    port map (
            O => \N__44857\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44854\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__10164\ : CascadeMux
    port map (
            O => \N__44851\,
            I => \N__44848\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44845\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44845\,
            I => \N__44841\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44837\
        );

    \I__10160\ : Span4Mux_h
    port map (
            O => \N__44841\,
            I => \N__44834\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44831\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44837\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__44834\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44831\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44821\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44821\,
            I => \N__44818\
        );

    \I__10153\ : Odrv12
    port map (
            O => \N__44818\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44815\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44808\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44805\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__44808\,
            I => \N__44799\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44799\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44804\,
            I => \N__44796\
        );

    \I__10146\ : Span4Mux_s3_v
    port map (
            O => \N__44799\,
            I => \N__44792\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44789\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44795\,
            I => \N__44786\
        );

    \I__10143\ : Span4Mux_h
    port map (
            O => \N__44792\,
            I => \N__44783\
        );

    \I__10142\ : Span4Mux_v
    port map (
            O => \N__44789\,
            I => \N__44778\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__44786\,
            I => \N__44778\
        );

    \I__10140\ : Sp12to4
    port map (
            O => \N__44783\,
            I => \N__44774\
        );

    \I__10139\ : Span4Mux_v
    port map (
            O => \N__44778\,
            I => \N__44771\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44777\,
            I => \N__44768\
        );

    \I__10137\ : Span12Mux_v
    port map (
            O => \N__44774\,
            I => \N__44765\
        );

    \I__10136\ : Sp12to4
    port map (
            O => \N__44771\,
            I => \N__44762\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44768\,
            I => \N__44759\
        );

    \I__10134\ : Span12Mux_v
    port map (
            O => \N__44765\,
            I => \N__44756\
        );

    \I__10133\ : Span12Mux_s7_h
    port map (
            O => \N__44762\,
            I => \N__44751\
        );

    \I__10132\ : Sp12to4
    port map (
            O => \N__44759\,
            I => \N__44751\
        );

    \I__10131\ : Span12Mux_h
    port map (
            O => \N__44756\,
            I => \N__44748\
        );

    \I__10130\ : Span12Mux_v
    port map (
            O => \N__44751\,
            I => \N__44745\
        );

    \I__10129\ : Odrv12
    port map (
            O => \N__44748\,
            I => start_stop_c
        );

    \I__10128\ : Odrv12
    port map (
            O => \N__44745\,
            I => start_stop_c
        );

    \I__10127\ : CascadeMux
    port map (
            O => \N__44740\,
            I => \N__44736\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44730\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44736\,
            I => \N__44725\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44735\,
            I => \N__44722\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44717\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44717\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44714\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44729\,
            I => \N__44708\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44728\,
            I => \N__44708\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44725\,
            I => \N__44705\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44722\,
            I => \N__44700\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__44717\,
            I => \N__44700\
        );

    \I__10115\ : Span4Mux_h
    port map (
            O => \N__44714\,
            I => \N__44697\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44713\,
            I => \N__44694\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44708\,
            I => phase_controller_inst1_state_4
        );

    \I__10112\ : Odrv12
    port map (
            O => \N__44705\,
            I => phase_controller_inst1_state_4
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__44700\,
            I => phase_controller_inst1_state_4
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__44697\,
            I => phase_controller_inst1_state_4
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44694\,
            I => phase_controller_inst1_state_4
        );

    \I__10108\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44679\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44682\,
            I => \N__44676\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__44679\,
            I => state_ns_i_a3_1
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__44676\,
            I => state_ns_i_a3_1
        );

    \I__10104\ : InMux
    port map (
            O => \N__44671\,
            I => \N__44667\
        );

    \I__10103\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44664\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44667\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44664\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44654\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44651\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44648\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44654\,
            I => \N__44643\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44651\,
            I => \N__44643\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44648\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__44643\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44638\,
            I => \N__44632\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44637\,
            I => \N__44632\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__44632\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44629\,
            I => \N__44626\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44626\,
            I => \N__44623\
        );

    \I__10088\ : Span4Mux_v
    port map (
            O => \N__44623\,
            I => \N__44620\
        );

    \I__10087\ : Span4Mux_h
    port map (
            O => \N__44620\,
            I => \N__44617\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__44617\,
            I => \N__44614\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__44614\,
            I => \pwm_generator_inst.O_0\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44608\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44608\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44602\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__44602\,
            I => \N__44599\
        );

    \I__10080\ : Span4Mux_v
    port map (
            O => \N__44599\,
            I => \N__44596\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__44596\,
            I => \N__44593\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__44593\,
            I => \N__44590\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__44590\,
            I => \pwm_generator_inst.O_1\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44587\,
            I => \N__44584\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44584\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44581\,
            I => \N__44578\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__44578\,
            I => \N__44575\
        );

    \I__10072\ : Span4Mux_h
    port map (
            O => \N__44575\,
            I => \N__44572\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__44572\,
            I => \N__44569\
        );

    \I__10070\ : Odrv4
    port map (
            O => \N__44569\,
            I => \pwm_generator_inst.O_2\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44563\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44563\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44560\,
            I => \N__44557\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44554\
        );

    \I__10065\ : Span12Mux_h
    port map (
            O => \N__44554\,
            I => \N__44551\
        );

    \I__10064\ : Odrv12
    port map (
            O => \N__44551\,
            I => \pwm_generator_inst.O_3\
        );

    \I__10063\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44545\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__44545\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__10061\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44539\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__44539\,
            I => \N__44536\
        );

    \I__10059\ : Span12Mux_s7_v
    port map (
            O => \N__44536\,
            I => \N__44533\
        );

    \I__10058\ : Odrv12
    port map (
            O => \N__44533\,
            I => \pwm_generator_inst.O_4\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44527\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__44527\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44524\,
            I => \N__44521\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44521\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__10053\ : CascadeMux
    port map (
            O => \N__44518\,
            I => \N__44515\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44512\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44506\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__44506\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__10048\ : CascadeMux
    port map (
            O => \N__44503\,
            I => \N__44500\
        );

    \I__10047\ : InMux
    port map (
            O => \N__44500\,
            I => \N__44497\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44497\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44494\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__44491\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__10043\ : IoInMux
    port map (
            O => \N__44488\,
            I => \N__44485\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__44485\,
            I => \N__44482\
        );

    \I__10041\ : Span4Mux_s3_v
    port map (
            O => \N__44482\,
            I => \N__44479\
        );

    \I__10040\ : Span4Mux_v
    port map (
            O => \N__44479\,
            I => \N__44476\
        );

    \I__10039\ : Span4Mux_v
    port map (
            O => \N__44476\,
            I => \N__44472\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44469\
        );

    \I__10037\ : Odrv4
    port map (
            O => \N__44472\,
            I => test_c
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44469\,
            I => test_c
        );

    \I__10035\ : CascadeMux
    port map (
            O => \N__44464\,
            I => \N__44461\
        );

    \I__10034\ : InMux
    port map (
            O => \N__44461\,
            I => \N__44458\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__44458\,
            I => \N__44455\
        );

    \I__10032\ : Odrv12
    port map (
            O => \N__44455\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44452\,
            I => \N__44449\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44449\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__10029\ : CascadeMux
    port map (
            O => \N__44446\,
            I => \N__44443\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44440\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__44440\,
            I => \N__44437\
        );

    \I__10026\ : Odrv12
    port map (
            O => \N__44437\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44431\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44431\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__44428\,
            I => \N__44425\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44425\,
            I => \N__44422\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44422\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44416\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__44416\,
            I => \N__44413\
        );

    \I__10018\ : Odrv12
    port map (
            O => \N__44413\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__10017\ : CascadeMux
    port map (
            O => \N__44410\,
            I => \N__44407\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44404\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__44404\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__10014\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44398\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44398\,
            I => \N__44395\
        );

    \I__10012\ : Odrv12
    port map (
            O => \N__44395\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__10011\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44389\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44386\
        );

    \I__10009\ : Odrv12
    port map (
            O => \N__44386\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__44383\,
            I => \N__44380\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44380\,
            I => \N__44377\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__44377\,
            I => \N__44374\
        );

    \I__10005\ : Odrv12
    port map (
            O => \N__44374\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44368\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44365\
        );

    \I__10002\ : Span4Mux_v
    port map (
            O => \N__44365\,
            I => \N__44362\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__44362\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__44359\,
            I => \N__44356\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44353\,
            I => \N__44350\
        );

    \I__9997\ : Odrv4
    port map (
            O => \N__44350\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__44347\,
            I => \N__44344\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44341\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44341\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44338\,
            I => \N__44335\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__44335\,
            I => \N__44332\
        );

    \I__9991\ : Odrv4
    port map (
            O => \N__44332\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__44329\,
            I => \N__44326\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44323\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44323\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44317\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__44317\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__44314\,
            I => \N__44311\
        );

    \I__9984\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44308\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__44308\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44302\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__44302\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__44299\,
            I => \N__44296\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44296\,
            I => \N__44293\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44290\
        );

    \I__9977\ : Odrv4
    port map (
            O => \N__44290\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44287\,
            I => \N__44284\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__44284\,
            I => \N__44281\
        );

    \I__9974\ : Odrv12
    port map (
            O => \N__44281\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__9973\ : CascadeMux
    port map (
            O => \N__44278\,
            I => \N__44275\
        );

    \I__9972\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44272\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__44272\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44266\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__44266\,
            I => \N__44263\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__44263\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__44260\,
            I => \N__44257\
        );

    \I__9966\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44254\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44254\,
            I => \N__44251\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__44251\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__9963\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44245\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44245\,
            I => \N__44242\
        );

    \I__9961\ : Span4Mux_v
    port map (
            O => \N__44242\,
            I => \N__44239\
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__44239\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__44236\,
            I => \N__44233\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44233\,
            I => \N__44230\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44230\,
            I => \N__44227\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__44227\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44224\,
            I => \N__44220\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44223\,
            I => \N__44217\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44212\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__44217\,
            I => \N__44209\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44204\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44215\,
            I => \N__44204\
        );

    \I__9949\ : Span4Mux_h
    port map (
            O => \N__44212\,
            I => \N__44201\
        );

    \I__9948\ : Span4Mux_h
    port map (
            O => \N__44209\,
            I => \N__44198\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__44204\,
            I => \N__44195\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__44201\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9945\ : Odrv4
    port map (
            O => \N__44198\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9944\ : Odrv12
    port map (
            O => \N__44195\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44183\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44180\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44186\,
            I => \N__44177\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44183\,
            I => \N__44172\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44180\,
            I => \N__44172\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__44177\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__9937\ : Odrv4
    port map (
            O => \N__44172\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44164\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44164\,
            I => \N__44160\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44156\
        );

    \I__9933\ : Span4Mux_v
    port map (
            O => \N__44160\,
            I => \N__44153\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44150\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44156\,
            I => \N__44147\
        );

    \I__9930\ : Span4Mux_h
    port map (
            O => \N__44153\,
            I => \N__44144\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44150\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__9928\ : Odrv12
    port map (
            O => \N__44147\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__44144\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__9926\ : CascadeMux
    port map (
            O => \N__44137\,
            I => \N__44132\
        );

    \I__9925\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44128\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44125\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44132\,
            I => \N__44122\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44131\,
            I => \N__44119\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__44128\,
            I => \N__44116\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__44125\,
            I => \N__44113\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__44122\,
            I => \N__44110\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44119\,
            I => \N__44101\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__44116\,
            I => \N__44101\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__44113\,
            I => \N__44101\
        );

    \I__9915\ : Span4Mux_v
    port map (
            O => \N__44110\,
            I => \N__44101\
        );

    \I__9914\ : Odrv4
    port map (
            O => \N__44101\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44098\,
            I => \N__44095\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44092\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__44092\,
            I => \N__44088\
        );

    \I__9910\ : InMux
    port map (
            O => \N__44091\,
            I => \N__44084\
        );

    \I__9909\ : Span4Mux_v
    port map (
            O => \N__44088\,
            I => \N__44081\
        );

    \I__9908\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44078\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__44084\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__9906\ : Odrv4
    port map (
            O => \N__44081\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44078\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__9904\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44066\
        );

    \I__9903\ : InMux
    port map (
            O => \N__44070\,
            I => \N__44062\
        );

    \I__9902\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44059\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__44066\,
            I => \N__44056\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44065\,
            I => \N__44053\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__44062\,
            I => \N__44050\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__44059\,
            I => \N__44047\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__44056\,
            I => \N__44042\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__44053\,
            I => \N__44042\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__44050\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__44047\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__44042\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__9892\ : InMux
    port map (
            O => \N__44035\,
            I => \N__44031\
        );

    \I__9891\ : InMux
    port map (
            O => \N__44034\,
            I => \N__44028\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__44031\,
            I => \N__44025\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__44021\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__44025\,
            I => \N__44018\
        );

    \I__9887\ : InMux
    port map (
            O => \N__44024\,
            I => \N__44015\
        );

    \I__9886\ : Span12Mux_h
    port map (
            O => \N__44021\,
            I => \N__44012\
        );

    \I__9885\ : Span4Mux_v
    port map (
            O => \N__44018\,
            I => \N__44009\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__44015\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__9883\ : Odrv12
    port map (
            O => \N__44012\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__44009\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__9881\ : InMux
    port map (
            O => \N__44002\,
            I => \N__43997\
        );

    \I__9880\ : InMux
    port map (
            O => \N__44001\,
            I => \N__43994\
        );

    \I__9879\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43991\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43987\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__43994\,
            I => \N__43984\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43991\,
            I => \N__43981\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43978\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__43987\,
            I => \N__43973\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__43984\,
            I => \N__43973\
        );

    \I__9872\ : Span4Mux_v
    port map (
            O => \N__43981\,
            I => \N__43970\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43978\,
            I => \N__43967\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__43973\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__43970\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__9868\ : Odrv4
    port map (
            O => \N__43967\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__9867\ : CascadeMux
    port map (
            O => \N__43960\,
            I => \N__43957\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43957\,
            I => \N__43954\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__43954\,
            I => \N__43951\
        );

    \I__9864\ : Span4Mux_v
    port map (
            O => \N__43951\,
            I => \N__43948\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__43948\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__9862\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43942\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43942\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__43939\,
            I => \N__43936\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43936\,
            I => \N__43933\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43930\
        );

    \I__9857\ : Odrv4
    port map (
            O => \N__43930\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43924\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43924\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43918\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__43918\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__9852\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43910\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43907\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43913\,
            I => \N__43904\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__43910\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__43907\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43904\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9846\ : CascadeMux
    port map (
            O => \N__43897\,
            I => \N__43892\
        );

    \I__9845\ : CascadeMux
    port map (
            O => \N__43896\,
            I => \N__43889\
        );

    \I__9844\ : CascadeMux
    port map (
            O => \N__43895\,
            I => \N__43885\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43892\,
            I => \N__43882\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43889\,
            I => \N__43879\
        );

    \I__9841\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43876\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43885\,
            I => \N__43873\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__43882\,
            I => \N__43864\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43879\,
            I => \N__43864\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__43876\,
            I => \N__43864\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43864\
        );

    \I__9835\ : Span4Mux_v
    port map (
            O => \N__43864\,
            I => \N__43861\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__43861\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9833\ : InMux
    port map (
            O => \N__43858\,
            I => \N__43854\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43850\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__43854\,
            I => \N__43847\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43843\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43850\,
            I => \N__43840\
        );

    \I__9828\ : Span4Mux_h
    port map (
            O => \N__43847\,
            I => \N__43837\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43834\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__43843\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__43840\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9824\ : Odrv4
    port map (
            O => \N__43837\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43834\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43822\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43818\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43814\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__43818\,
            I => \N__43811\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43808\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43814\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__43811\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43808\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43796\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43793\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43790\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__43796\,
            I => \N__43785\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43793\,
            I => \N__43785\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43790\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__9808\ : Odrv12
    port map (
            O => \N__43785\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43780\,
            I => \N__43776\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43773\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43776\,
            I => \N__43768\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43773\,
            I => \N__43765\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43772\,
            I => \N__43762\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43771\,
            I => \N__43759\
        );

    \I__9801\ : Span4Mux_h
    port map (
            O => \N__43768\,
            I => \N__43754\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__43765\,
            I => \N__43754\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43762\,
            I => \N__43751\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43759\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__9797\ : Odrv4
    port map (
            O => \N__43754\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__9796\ : Odrv12
    port map (
            O => \N__43751\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43740\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43736\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43740\,
            I => \N__43733\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43739\,
            I => \N__43730\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__43736\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9790\ : Odrv4
    port map (
            O => \N__43733\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43730\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9788\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43718\
        );

    \I__9787\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43715\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43712\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__43718\,
            I => \N__43707\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43707\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43712\,
            I => \N__43703\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__43707\,
            I => \N__43700\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43706\,
            I => \N__43697\
        );

    \I__9780\ : Odrv4
    port map (
            O => \N__43703\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9779\ : Odrv4
    port map (
            O => \N__43700\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__43697\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43686\
        );

    \I__9776\ : InMux
    port map (
            O => \N__43689\,
            I => \N__43682\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43686\,
            I => \N__43679\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43676\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43682\,
            I => \N__43671\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__43679\,
            I => \N__43671\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43668\
        );

    \I__9770\ : Odrv4
    port map (
            O => \N__43671\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__9769\ : Odrv4
    port map (
            O => \N__43668\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43657\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43654\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43651\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43648\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43657\,
            I => \N__43643\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43654\,
            I => \N__43643\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43651\,
            I => \N__43638\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__43648\,
            I => \N__43638\
        );

    \I__9760\ : Span4Mux_v
    port map (
            O => \N__43643\,
            I => \N__43635\
        );

    \I__9759\ : Span4Mux_v
    port map (
            O => \N__43638\,
            I => \N__43632\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__43635\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9757\ : Odrv4
    port map (
            O => \N__43632\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43621\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43621\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__43621\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__9753\ : CascadeMux
    port map (
            O => \N__43618\,
            I => \N__43615\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43615\,
            I => \N__43609\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43614\,
            I => \N__43609\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__43609\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43602\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43605\,
            I => \N__43599\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43602\,
            I => \N__43592\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43599\,
            I => \N__43592\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43598\,
            I => \N__43589\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43597\,
            I => \N__43586\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__43592\,
            I => \N__43583\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43589\,
            I => \N__43580\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__43586\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__43583\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__9739\ : Odrv12
    port map (
            O => \N__43580\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43569\
        );

    \I__9737\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43566\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43569\,
            I => \N__43559\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43559\
        );

    \I__9734\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43556\
        );

    \I__9733\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43553\
        );

    \I__9732\ : Span4Mux_v
    port map (
            O => \N__43559\,
            I => \N__43550\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__43556\,
            I => \N__43547\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43553\,
            I => \N__43544\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__43550\,
            I => \N__43539\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__43547\,
            I => \N__43539\
        );

    \I__9727\ : Odrv4
    port map (
            O => \N__43544\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9726\ : Odrv4
    port map (
            O => \N__43539\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__43534\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\
        );

    \I__9724\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43528\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__43528\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__9722\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43522\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__43522\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__43519\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43513\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__43513\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__43510\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__9716\ : InMux
    port map (
            O => \N__43507\,
            I => \N__43502\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43506\,
            I => \N__43499\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43505\,
            I => \N__43496\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__43502\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43499\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43496\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43485\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43482\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43485\,
            I => \N__43476\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__43482\,
            I => \N__43476\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43481\,
            I => \N__43473\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__43476\,
            I => \N__43467\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__43473\,
            I => \N__43467\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43464\
        );

    \I__9702\ : Span4Mux_h
    port map (
            O => \N__43467\,
            I => \N__43461\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43458\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__43461\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9699\ : Odrv12
    port map (
            O => \N__43458\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9698\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43450\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__43450\,
            I => \N__43445\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43442\
        );

    \I__9695\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43439\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__43445\,
            I => \N__43436\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__43442\,
            I => \N__43433\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__43439\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__43436\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__9690\ : Odrv12
    port map (
            O => \N__43433\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__9689\ : InMux
    port map (
            O => \N__43426\,
            I => \N__43423\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__43423\,
            I => \N__43419\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43422\,
            I => \N__43416\
        );

    \I__9686\ : Span4Mux_v
    port map (
            O => \N__43419\,
            I => \N__43409\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43416\,
            I => \N__43409\
        );

    \I__9684\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43406\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43414\,
            I => \N__43403\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__43409\,
            I => \N__43398\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43398\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43403\,
            I => \N__43395\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__43398\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__9678\ : Odrv12
    port map (
            O => \N__43395\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__43390\,
            I => \N__43387\
        );

    \I__9676\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43384\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43381\
        );

    \I__9674\ : Span4Mux_v
    port map (
            O => \N__43381\,
            I => \N__43378\
        );

    \I__9673\ : Sp12to4
    port map (
            O => \N__43378\,
            I => \N__43375\
        );

    \I__9672\ : Span12Mux_h
    port map (
            O => \N__43375\,
            I => \N__43372\
        );

    \I__9671\ : Odrv12
    port map (
            O => \N__43372\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__9670\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43366\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__43366\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__9668\ : InMux
    port map (
            O => \N__43363\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43360\,
            I => \N__43357\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__43357\,
            I => \N__43354\
        );

    \I__9665\ : Span4Mux_v
    port map (
            O => \N__43354\,
            I => \N__43351\
        );

    \I__9664\ : Sp12to4
    port map (
            O => \N__43351\,
            I => \N__43348\
        );

    \I__9663\ : Span12Mux_h
    port map (
            O => \N__43348\,
            I => \N__43345\
        );

    \I__9662\ : Odrv12
    port map (
            O => \N__43345\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__43342\,
            I => \N__43336\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__43341\,
            I => \N__43332\
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__43340\,
            I => \N__43328\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43324\
        );

    \I__9657\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43311\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43311\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43311\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43331\,
            I => \N__43311\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43328\,
            I => \N__43311\
        );

    \I__9652\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43311\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__43324\,
            I => \N__43308\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N__43304\
        );

    \I__9649\ : Span12Mux_s7_v
    port map (
            O => \N__43308\,
            I => \N__43301\
        );

    \I__9648\ : InMux
    port map (
            O => \N__43307\,
            I => \N__43298\
        );

    \I__9647\ : Span4Mux_h
    port map (
            O => \N__43304\,
            I => \N__43295\
        );

    \I__9646\ : Span12Mux_h
    port map (
            O => \N__43301\,
            I => \N__43290\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__43298\,
            I => \N__43290\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__43295\,
            I => \N__43287\
        );

    \I__9643\ : Span12Mux_h
    port map (
            O => \N__43290\,
            I => \N__43284\
        );

    \I__9642\ : Span4Mux_h
    port map (
            O => \N__43287\,
            I => \N__43281\
        );

    \I__9641\ : Odrv12
    port map (
            O => \N__43284\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__43281\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__9639\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43273\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__43273\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__9637\ : InMux
    port map (
            O => \N__43270\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43267\,
            I => \N__43264\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__43264\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43258\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43258\,
            I => \N__43255\
        );

    \I__9632\ : Span4Mux_v
    port map (
            O => \N__43255\,
            I => \N__43252\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__43252\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43249\,
            I => \bfn_16_29_0_\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43246\,
            I => \N__43243\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43239\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43236\
        );

    \I__9626\ : Odrv4
    port map (
            O => \N__43239\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__43236\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__9624\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43228\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__43228\,
            I => \N__43225\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__43225\,
            I => \N__43222\
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__43222\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43216\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__43216\,
            I => \N__43213\
        );

    \I__9618\ : Span4Mux_v
    port map (
            O => \N__43213\,
            I => \N__43210\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__43210\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43207\,
            I => \N__43202\
        );

    \I__9615\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43199\
        );

    \I__9614\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43196\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43202\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__43199\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__43196\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__9610\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43184\
        );

    \I__9609\ : InMux
    port map (
            O => \N__43188\,
            I => \N__43181\
        );

    \I__9608\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43178\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__43184\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__43181\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__43178\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43171\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43168\,
            I => \N__43165\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__43165\,
            I => \N__43162\
        );

    \I__9601\ : Span4Mux_v
    port map (
            O => \N__43162\,
            I => \N__43159\
        );

    \I__9600\ : Sp12to4
    port map (
            O => \N__43159\,
            I => \N__43156\
        );

    \I__9599\ : Odrv12
    port map (
            O => \N__43156\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__43153\,
            I => \N__43150\
        );

    \I__9597\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43147\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__43147\,
            I => \N__43144\
        );

    \I__9595\ : Span4Mux_v
    port map (
            O => \N__43144\,
            I => \N__43141\
        );

    \I__9594\ : Sp12to4
    port map (
            O => \N__43141\,
            I => \N__43138\
        );

    \I__9593\ : Span12Mux_h
    port map (
            O => \N__43138\,
            I => \N__43135\
        );

    \I__9592\ : Odrv12
    port map (
            O => \N__43135\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__9591\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43129\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43129\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__9589\ : InMux
    port map (
            O => \N__43126\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43123\,
            I => \N__43120\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__43120\,
            I => \N__43117\
        );

    \I__9586\ : Span4Mux_v
    port map (
            O => \N__43117\,
            I => \N__43114\
        );

    \I__9585\ : Sp12to4
    port map (
            O => \N__43114\,
            I => \N__43111\
        );

    \I__9584\ : Odrv12
    port map (
            O => \N__43111\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__43108\,
            I => \N__43105\
        );

    \I__9582\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43102\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43102\,
            I => \N__43099\
        );

    \I__9580\ : Span4Mux_v
    port map (
            O => \N__43099\,
            I => \N__43096\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__43096\,
            I => \N__43093\
        );

    \I__9578\ : Span4Mux_h
    port map (
            O => \N__43093\,
            I => \N__43090\
        );

    \I__9577\ : Span4Mux_h
    port map (
            O => \N__43090\,
            I => \N__43087\
        );

    \I__9576\ : Odrv4
    port map (
            O => \N__43087\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__9575\ : InMux
    port map (
            O => \N__43084\,
            I => \N__43081\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43081\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__9573\ : InMux
    port map (
            O => \N__43078\,
            I => \bfn_16_28_0_\
        );

    \I__9572\ : InMux
    port map (
            O => \N__43075\,
            I => \N__43072\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__43072\,
            I => \N__43069\
        );

    \I__9570\ : Span4Mux_h
    port map (
            O => \N__43069\,
            I => \N__43066\
        );

    \I__9569\ : Span4Mux_h
    port map (
            O => \N__43066\,
            I => \N__43063\
        );

    \I__9568\ : Span4Mux_h
    port map (
            O => \N__43063\,
            I => \N__43060\
        );

    \I__9567\ : Odrv4
    port map (
            O => \N__43060\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__9566\ : CascadeMux
    port map (
            O => \N__43057\,
            I => \N__43054\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43051\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43051\,
            I => \N__43048\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__43048\,
            I => \N__43045\
        );

    \I__9562\ : Sp12to4
    port map (
            O => \N__43045\,
            I => \N__43042\
        );

    \I__9561\ : Span12Mux_h
    port map (
            O => \N__43042\,
            I => \N__43039\
        );

    \I__9560\ : Odrv12
    port map (
            O => \N__43039\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43036\,
            I => \N__43033\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__43033\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__9557\ : InMux
    port map (
            O => \N__43030\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__9556\ : CascadeMux
    port map (
            O => \N__43027\,
            I => \N__43024\
        );

    \I__9555\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43021\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43021\,
            I => \N__43018\
        );

    \I__9553\ : Span4Mux_v
    port map (
            O => \N__43018\,
            I => \N__43015\
        );

    \I__9552\ : Span4Mux_h
    port map (
            O => \N__43015\,
            I => \N__43012\
        );

    \I__9551\ : Span4Mux_h
    port map (
            O => \N__43012\,
            I => \N__43009\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__43006\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__9548\ : InMux
    port map (
            O => \N__43003\,
            I => \N__43000\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__43000\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42997\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42991\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42991\,
            I => \N__42988\
        );

    \I__9543\ : Span4Mux_v
    port map (
            O => \N__42988\,
            I => \N__42985\
        );

    \I__9542\ : Sp12to4
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__9541\ : Span12Mux_h
    port map (
            O => \N__42982\,
            I => \N__42979\
        );

    \I__9540\ : Odrv12
    port map (
            O => \N__42979\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42973\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42973\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__9537\ : InMux
    port map (
            O => \N__42970\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42961\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__42961\,
            I => \N__42958\
        );

    \I__9533\ : Span12Mux_s6_v
    port map (
            O => \N__42958\,
            I => \N__42955\
        );

    \I__9532\ : Span12Mux_h
    port map (
            O => \N__42955\,
            I => \N__42952\
        );

    \I__9531\ : Odrv12
    port map (
            O => \N__42952\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42946\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42946\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__9528\ : InMux
    port map (
            O => \N__42943\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42937\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__42937\,
            I => \N__42934\
        );

    \I__9525\ : Span4Mux_h
    port map (
            O => \N__42934\,
            I => \N__42931\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__42931\,
            I => \N__42928\
        );

    \I__9523\ : Sp12to4
    port map (
            O => \N__42928\,
            I => \N__42925\
        );

    \I__9522\ : Odrv12
    port map (
            O => \N__42925\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42919\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__42919\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42916\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__42913\,
            I => \N__42910\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42906\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42903\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__42906\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__42903\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42895\,
            I => \N__42892\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__42892\,
            I => \N__42889\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__42889\,
            I => \N__42886\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__42886\,
            I => \N__42883\
        );

    \I__9508\ : Span4Mux_h
    port map (
            O => \N__42883\,
            I => \N__42880\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__42880\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__9506\ : CascadeMux
    port map (
            O => \N__42877\,
            I => \N__42874\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42868\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__42868\,
            I => \N__42865\
        );

    \I__9502\ : Span4Mux_h
    port map (
            O => \N__42865\,
            I => \N__42862\
        );

    \I__9501\ : Span4Mux_h
    port map (
            O => \N__42862\,
            I => \N__42859\
        );

    \I__9500\ : Odrv4
    port map (
            O => \N__42859\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42853\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42853\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42847\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42844\
        );

    \I__9495\ : Span4Mux_h
    port map (
            O => \N__42844\,
            I => \N__42841\
        );

    \I__9494\ : Span4Mux_h
    port map (
            O => \N__42841\,
            I => \N__42838\
        );

    \I__9493\ : Span4Mux_h
    port map (
            O => \N__42838\,
            I => \N__42835\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__42835\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__42832\,
            I => \N__42829\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42829\,
            I => \N__42826\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42826\,
            I => \N__42823\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__42823\,
            I => \N__42820\
        );

    \I__9487\ : Sp12to4
    port map (
            O => \N__42820\,
            I => \N__42817\
        );

    \I__9486\ : Span12Mux_h
    port map (
            O => \N__42817\,
            I => \N__42814\
        );

    \I__9485\ : Odrv12
    port map (
            O => \N__42814\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__42811\,
            I => \N__42808\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42805\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__42805\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42802\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42796\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__42796\,
            I => \N__42793\
        );

    \I__9478\ : Span4Mux_v
    port map (
            O => \N__42793\,
            I => \N__42790\
        );

    \I__9477\ : Sp12to4
    port map (
            O => \N__42790\,
            I => \N__42787\
        );

    \I__9476\ : Span12Mux_h
    port map (
            O => \N__42787\,
            I => \N__42784\
        );

    \I__9475\ : Odrv12
    port map (
            O => \N__42784\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__9474\ : CascadeMux
    port map (
            O => \N__42781\,
            I => \N__42778\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42775\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42775\,
            I => \N__42772\
        );

    \I__9471\ : Span4Mux_h
    port map (
            O => \N__42772\,
            I => \N__42769\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__42769\,
            I => \N__42766\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__42766\,
            I => \N__42763\
        );

    \I__9468\ : Odrv4
    port map (
            O => \N__42763\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42760\,
            I => \N__42757\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__42757\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__9465\ : InMux
    port map (
            O => \N__42754\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42751\,
            I => \N__42748\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42748\,
            I => \N__42745\
        );

    \I__9462\ : Span4Mux_v
    port map (
            O => \N__42745\,
            I => \N__42742\
        );

    \I__9461\ : Sp12to4
    port map (
            O => \N__42742\,
            I => \N__42739\
        );

    \I__9460\ : Span12Mux_h
    port map (
            O => \N__42739\,
            I => \N__42736\
        );

    \I__9459\ : Odrv12
    port map (
            O => \N__42736\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__42733\,
            I => \N__42730\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42730\,
            I => \N__42727\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42727\,
            I => \N__42724\
        );

    \I__9455\ : Span12Mux_h
    port map (
            O => \N__42724\,
            I => \N__42721\
        );

    \I__9454\ : Odrv12
    port map (
            O => \N__42721\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__9453\ : CascadeMux
    port map (
            O => \N__42718\,
            I => \N__42715\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42712\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42712\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42709\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42703\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42703\,
            I => \N__42700\
        );

    \I__9447\ : Span12Mux_s7_v
    port map (
            O => \N__42700\,
            I => \N__42697\
        );

    \I__9446\ : Span12Mux_h
    port map (
            O => \N__42697\,
            I => \N__42694\
        );

    \I__9445\ : Odrv12
    port map (
            O => \N__42694\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__9444\ : CascadeMux
    port map (
            O => \N__42691\,
            I => \N__42688\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42688\,
            I => \N__42685\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42685\,
            I => \N__42682\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__42682\,
            I => \N__42679\
        );

    \I__9440\ : Span4Mux_h
    port map (
            O => \N__42679\,
            I => \N__42676\
        );

    \I__9439\ : Span4Mux_h
    port map (
            O => \N__42676\,
            I => \N__42673\
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__42673\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42667\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42667\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42664\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42661\,
            I => \N__42658\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42655\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__42655\,
            I => \N__42652\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__42652\,
            I => \N__42649\
        );

    \I__9430\ : Sp12to4
    port map (
            O => \N__42649\,
            I => \N__42646\
        );

    \I__9429\ : Odrv12
    port map (
            O => \N__42646\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__42643\,
            I => \N__42640\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42637\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42634\
        );

    \I__9425\ : Span4Mux_v
    port map (
            O => \N__42634\,
            I => \N__42631\
        );

    \I__9424\ : Sp12to4
    port map (
            O => \N__42631\,
            I => \N__42628\
        );

    \I__9423\ : Odrv12
    port map (
            O => \N__42628\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42622\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42622\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42619\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42613\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42613\,
            I => \N__42610\
        );

    \I__9417\ : Span12Mux_s5_v
    port map (
            O => \N__42610\,
            I => \N__42607\
        );

    \I__9416\ : Odrv12
    port map (
            O => \N__42607\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__9415\ : CascadeMux
    port map (
            O => \N__42604\,
            I => \N__42601\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42598\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42595\
        );

    \I__9412\ : Span4Mux_v
    port map (
            O => \N__42595\,
            I => \N__42592\
        );

    \I__9411\ : Sp12to4
    port map (
            O => \N__42592\,
            I => \N__42589\
        );

    \I__9410\ : Span12Mux_h
    port map (
            O => \N__42589\,
            I => \N__42586\
        );

    \I__9409\ : Odrv12
    port map (
            O => \N__42586\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42580\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42580\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__9406\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42574\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__42574\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__9404\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42568\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__42568\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__9402\ : CascadeMux
    port map (
            O => \N__42565\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\
        );

    \I__9401\ : InMux
    port map (
            O => \N__42562\,
            I => \N__42559\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__42559\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__9399\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42551\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42548\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42545\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42551\,
            I => \N__42538\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42548\,
            I => \N__42538\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__42545\,
            I => \N__42538\
        );

    \I__9393\ : Span4Mux_v
    port map (
            O => \N__42538\,
            I => \N__42535\
        );

    \I__9392\ : Sp12to4
    port map (
            O => \N__42535\,
            I => \N__42532\
        );

    \I__9391\ : Span12Mux_h
    port map (
            O => \N__42532\,
            I => \N__42529\
        );

    \I__9390\ : Span12Mux_v
    port map (
            O => \N__42529\,
            I => \N__42526\
        );

    \I__9389\ : Odrv12
    port map (
            O => \N__42526\,
            I => il_min_comp2_c
        );

    \I__9388\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42520\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__42520\,
            I => \N__42517\
        );

    \I__9386\ : Span4Mux_v
    port map (
            O => \N__42517\,
            I => \N__42513\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42510\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__42513\,
            I => \N__42505\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42510\,
            I => \N__42505\
        );

    \I__9382\ : Odrv4
    port map (
            O => \N__42505\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__9381\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42498\
        );

    \I__9380\ : CascadeMux
    port map (
            O => \N__42501\,
            I => \N__42495\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__9378\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42488\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__42492\,
            I => \N__42485\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42491\,
            I => \N__42481\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__42488\,
            I => \N__42478\
        );

    \I__9374\ : Span4Mux_v
    port map (
            O => \N__42485\,
            I => \N__42475\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42484\,
            I => \N__42472\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__42481\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__42478\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__42475\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__42472\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42463\,
            I => \N__42458\
        );

    \I__9367\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42455\
        );

    \I__9366\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42452\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42458\,
            I => \N__42449\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42455\,
            I => \N__42444\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__42452\,
            I => \N__42444\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__42449\,
            I => \N__42440\
        );

    \I__9361\ : Span4Mux_v
    port map (
            O => \N__42444\,
            I => \N__42437\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42432\
        );

    \I__9359\ : Sp12to4
    port map (
            O => \N__42440\,
            I => \N__42427\
        );

    \I__9358\ : Sp12to4
    port map (
            O => \N__42437\,
            I => \N__42427\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42436\,
            I => \N__42424\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42435\,
            I => \N__42420\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__42432\,
            I => \N__42417\
        );

    \I__9354\ : Span12Mux_h
    port map (
            O => \N__42427\,
            I => \N__42412\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__42424\,
            I => \N__42412\
        );

    \I__9352\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42409\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__42420\,
            I => state_3
        );

    \I__9350\ : Odrv4
    port map (
            O => \N__42417\,
            I => state_3
        );

    \I__9349\ : Odrv12
    port map (
            O => \N__42412\,
            I => state_3
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42409\,
            I => state_3
        );

    \I__9347\ : IoInMux
    port map (
            O => \N__42400\,
            I => \N__42397\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__42397\,
            I => \N__42394\
        );

    \I__9345\ : Span4Mux_s1_v
    port map (
            O => \N__42394\,
            I => \N__42391\
        );

    \I__9344\ : Span4Mux_v
    port map (
            O => \N__42391\,
            I => \N__42388\
        );

    \I__9343\ : Span4Mux_v
    port map (
            O => \N__42388\,
            I => \N__42384\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42381\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__42384\,
            I => test22_c
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__42381\,
            I => test22_c
        );

    \I__9339\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42348\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42331\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42331\
        );

    \I__9336\ : InMux
    port map (
            O => \N__42373\,
            I => \N__42331\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42372\,
            I => \N__42331\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42331\
        );

    \I__9333\ : InMux
    port map (
            O => \N__42370\,
            I => \N__42331\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42331\
        );

    \I__9331\ : InMux
    port map (
            O => \N__42368\,
            I => \N__42331\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42316\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42316\
        );

    \I__9328\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42316\
        );

    \I__9327\ : InMux
    port map (
            O => \N__42364\,
            I => \N__42316\
        );

    \I__9326\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42316\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42362\,
            I => \N__42316\
        );

    \I__9324\ : InMux
    port map (
            O => \N__42361\,
            I => \N__42316\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__42360\,
            I => \N__42313\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__42359\,
            I => \N__42306\
        );

    \I__9321\ : CascadeMux
    port map (
            O => \N__42358\,
            I => \N__42302\
        );

    \I__9320\ : CascadeMux
    port map (
            O => \N__42357\,
            I => \N__42299\
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__42356\,
            I => \N__42296\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42355\,
            I => \N__42291\
        );

    \I__9317\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42291\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42284\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42352\,
            I => \N__42284\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42284\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42348\,
            I => \N__42277\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42277\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__42316\,
            I => \N__42277\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42313\,
            I => \N__42274\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42271\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42256\
        );

    \I__9307\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42256\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42309\,
            I => \N__42256\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42256\
        );

    \I__9304\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42256\
        );

    \I__9303\ : InMux
    port map (
            O => \N__42302\,
            I => \N__42256\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42299\,
            I => \N__42256\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42253\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42247\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42284\,
            I => \N__42247\
        );

    \I__9298\ : Span4Mux_v
    port map (
            O => \N__42277\,
            I => \N__42244\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__42274\,
            I => \N__42239\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42271\,
            I => \N__42239\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42256\,
            I => \N__42236\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42233\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__42252\,
            I => \N__42230\
        );

    \I__9292\ : Span4Mux_v
    port map (
            O => \N__42247\,
            I => \N__42227\
        );

    \I__9291\ : Sp12to4
    port map (
            O => \N__42244\,
            I => \N__42224\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__42239\,
            I => \N__42221\
        );

    \I__9289\ : Span4Mux_h
    port map (
            O => \N__42236\,
            I => \N__42218\
        );

    \I__9288\ : Span4Mux_h
    port map (
            O => \N__42233\,
            I => \N__42215\
        );

    \I__9287\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42212\
        );

    \I__9286\ : Sp12to4
    port map (
            O => \N__42227\,
            I => \N__42209\
        );

    \I__9285\ : Span12Mux_s8_h
    port map (
            O => \N__42224\,
            I => \N__42206\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__42221\,
            I => \N_19_1\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__42218\,
            I => \N_19_1\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__42215\,
            I => \N_19_1\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42212\,
            I => \N_19_1\
        );

    \I__9280\ : Odrv12
    port map (
            O => \N__42209\,
            I => \N_19_1\
        );

    \I__9279\ : Odrv12
    port map (
            O => \N__42206\,
            I => \N_19_1\
        );

    \I__9278\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42189\
        );

    \I__9277\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42186\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__42189\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__42186\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__9274\ : InMux
    port map (
            O => \N__42181\,
            I => \N__42175\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42175\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__42175\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__42172\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42166\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42163\
        );

    \I__9268\ : Odrv12
    port map (
            O => \N__42163\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__9267\ : InMux
    port map (
            O => \N__42160\,
            I => \N__42156\
        );

    \I__9266\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42153\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__42156\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__42153\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__9263\ : InMux
    port map (
            O => \N__42148\,
            I => \N__42141\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42141\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42137\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42141\,
            I => \N__42134\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42131\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__42137\,
            I => \N__42128\
        );

    \I__9257\ : Span4Mux_h
    port map (
            O => \N__42134\,
            I => \N__42125\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42131\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__9255\ : Odrv12
    port map (
            O => \N__42128\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__42125\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__9253\ : CascadeMux
    port map (
            O => \N__42118\,
            I => \N__42115\
        );

    \I__9252\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42112\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42112\,
            I => \N__42108\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42111\,
            I => \N__42105\
        );

    \I__9249\ : Odrv4
    port map (
            O => \N__42108\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__42105\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42100\,
            I => \N__42097\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__42097\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__9245\ : CascadeMux
    port map (
            O => \N__42094\,
            I => \N__42090\
        );

    \I__9244\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42087\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42082\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42087\,
            I => \N__42079\
        );

    \I__9241\ : InMux
    port map (
            O => \N__42086\,
            I => \N__42074\
        );

    \I__9240\ : InMux
    port map (
            O => \N__42085\,
            I => \N__42074\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__42082\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__42079\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__42074\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__42067\,
            I => \N__42064\
        );

    \I__9235\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42061\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42061\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__9233\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42055\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__42055\,
            I => \N__42052\
        );

    \I__9231\ : Span4Mux_h
    port map (
            O => \N__42052\,
            I => \N__42049\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__42049\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42046\,
            I => \N__42042\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42039\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__42042\,
            I => \N__42034\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__42034\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__42034\,
            I => \N__42030\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42027\
        );

    \I__9223\ : Sp12to4
    port map (
            O => \N__42030\,
            I => \N__42022\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__42022\
        );

    \I__9221\ : Span12Mux_h
    port map (
            O => \N__42022\,
            I => \N__42019\
        );

    \I__9220\ : Span12Mux_v
    port map (
            O => \N__42019\,
            I => \N__42016\
        );

    \I__9219\ : Odrv12
    port map (
            O => \N__42016\,
            I => il_max_comp2_c
        );

    \I__9218\ : InMux
    port map (
            O => \N__42013\,
            I => \N__42010\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__42010\,
            I => \N__42006\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__42009\,
            I => \N__42002\
        );

    \I__9215\ : Span4Mux_v
    port map (
            O => \N__42006\,
            I => \N__41999\
        );

    \I__9214\ : CascadeMux
    port map (
            O => \N__42005\,
            I => \N__41996\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41993\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__41999\,
            I => \N__41990\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41986\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41993\,
            I => \N__41981\
        );

    \I__9209\ : Span4Mux_v
    port map (
            O => \N__41990\,
            I => \N__41981\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41978\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41986\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9206\ : Odrv4
    port map (
            O => \N__41981\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41978\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41971\,
            I => \N__41968\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__41968\,
            I => \N__41964\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41961\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__41964\,
            I => \N__41958\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41961\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__41958\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41950\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41950\,
            I => \N__41946\
        );

    \I__9196\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41943\
        );

    \I__9195\ : Odrv4
    port map (
            O => \N__41946\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41943\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__9193\ : CascadeMux
    port map (
            O => \N__41938\,
            I => \N__41935\
        );

    \I__9192\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41932\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__41932\,
            I => \N__41928\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41925\
        );

    \I__9189\ : Odrv4
    port map (
            O => \N__41928\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41925\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41910\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41907\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__41910\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41907\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41899\,
            I => \N__41895\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41898\,
            I => \N__41892\
        );

    \I__9178\ : Span4Mux_v
    port map (
            O => \N__41895\,
            I => \N__41889\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41892\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9176\ : Odrv4
    port map (
            O => \N__41889\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41881\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41881\,
            I => \N__41875\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41870\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41870\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41878\,
            I => \N__41867\
        );

    \I__9170\ : Span4Mux_h
    port map (
            O => \N__41875\,
            I => \N__41862\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__41870\,
            I => \N__41862\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__41867\,
            I => \N__41859\
        );

    \I__9167\ : Odrv4
    port map (
            O => \N__41862\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__41859\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9165\ : CascadeMux
    port map (
            O => \N__41854\,
            I => \N__41851\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41845\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41845\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41845\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41842\,
            I => \N__41838\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41835\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__41838\,
            I => \N__41831\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41828\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41825\
        );

    \I__9156\ : Odrv12
    port map (
            O => \N__41831\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__41828\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41825\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__41818\,
            I => \N__41815\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41811\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41808\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__41811\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__41808\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9148\ : CascadeMux
    port map (
            O => \N__41803\,
            I => \N__41798\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41802\,
            I => \N__41795\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41790\
        );

    \I__9145\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41787\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__41795\,
            I => \N__41784\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41794\,
            I => \N__41779\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41779\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41790\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41787\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9139\ : Odrv4
    port map (
            O => \N__41784\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41779\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41767\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41767\,
            I => \N__41762\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41766\,
            I => \N__41755\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41755\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__41762\,
            I => \N__41752\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41749\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41746\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41755\,
            I => \N__41743\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__41752\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41749\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__41746\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9126\ : Odrv12
    port map (
            O => \N__41743\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41731\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41727\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41724\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__41727\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41724\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41719\,
            I => \N__41714\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41711\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41717\,
            I => \N__41708\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41714\,
            I => \N__41705\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41711\,
            I => \N__41700\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41708\,
            I => \N__41700\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__41705\,
            I => \N__41697\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__41700\,
            I => \N__41694\
        );

    \I__9112\ : Sp12to4
    port map (
            O => \N__41697\,
            I => \N__41689\
        );

    \I__9111\ : Sp12to4
    port map (
            O => \N__41694\,
            I => \N__41689\
        );

    \I__9110\ : Span12Mux_h
    port map (
            O => \N__41689\,
            I => \N__41686\
        );

    \I__9109\ : Span12Mux_v
    port map (
            O => \N__41686\,
            I => \N__41683\
        );

    \I__9108\ : Odrv12
    port map (
            O => \N__41683\,
            I => il_max_comp1_c
        );

    \I__9107\ : InMux
    port map (
            O => \N__41680\,
            I => \N__41673\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41673\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41670\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41673\,
            I => \N__41665\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__41670\,
            I => \N__41665\
        );

    \I__9102\ : Span4Mux_v
    port map (
            O => \N__41665\,
            I => \N__41662\
        );

    \I__9101\ : Sp12to4
    port map (
            O => \N__41662\,
            I => \N__41659\
        );

    \I__9100\ : Span12Mux_h
    port map (
            O => \N__41659\,
            I => \N__41656\
        );

    \I__9099\ : Span12Mux_v
    port map (
            O => \N__41656\,
            I => \N__41653\
        );

    \I__9098\ : Odrv12
    port map (
            O => \N__41653\,
            I => il_min_comp1_c
        );

    \I__9097\ : CascadeMux
    port map (
            O => \N__41650\,
            I => \N__41647\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41643\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41639\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41636\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41633\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__41639\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__41636\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__41633\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41623\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41623\,
            I => \N__41620\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__41620\,
            I => \N__41614\
        );

    \I__9086\ : InMux
    port map (
            O => \N__41619\,
            I => \N__41609\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41618\,
            I => \N__41609\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41606\
        );

    \I__9083\ : Odrv4
    port map (
            O => \N__41614\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41609\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__41606\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41595\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41592\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41595\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__41592\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41584\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41584\,
            I => \N__41579\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41573\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41573\
        );

    \I__9072\ : Span4Mux_v
    port map (
            O => \N__41579\,
            I => \N__41570\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41567\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41564\
        );

    \I__9069\ : Odrv4
    port map (
            O => \N__41570\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__41567\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__41564\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41554\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__41554\,
            I => \N__41550\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41547\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__41550\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__41547\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__41542\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41539\,
            I => \N__41534\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41531\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41528\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__41534\,
            I => \N__41523\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__41531\,
            I => \N__41523\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41528\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9054\ : Odrv12
    port map (
            O => \N__41523\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41513\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41517\,
            I => \N__41510\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41516\,
            I => \N__41507\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41513\,
            I => \N__41504\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__41510\,
            I => \N__41501\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__41507\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__9047\ : Odrv4
    port map (
            O => \N__41504\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__41501\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41490\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41486\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41482\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41479\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41486\,
            I => \N__41476\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41473\
        );

    \I__9039\ : Span4Mux_v
    port map (
            O => \N__41482\,
            I => \N__41470\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41465\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__41476\,
            I => \N__41465\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41462\
        );

    \I__9035\ : Odrv4
    port map (
            O => \N__41470\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9034\ : Odrv4
    port map (
            O => \N__41465\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__41462\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41449\
        );

    \I__9031\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41449\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41449\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41446\,
            I => \N__41441\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41438\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41435\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41441\,
            I => \N__41432\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41438\,
            I => \N__41428\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__41435\,
            I => \N__41425\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__41432\,
            I => \N__41422\
        );

    \I__9022\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41419\
        );

    \I__9021\ : Span4Mux_h
    port map (
            O => \N__41428\,
            I => \N__41414\
        );

    \I__9020\ : Span4Mux_h
    port map (
            O => \N__41425\,
            I => \N__41414\
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__41422\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41419\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__41414\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41402\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41399\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41396\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41402\,
            I => \N__41393\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__41399\,
            I => \N__41390\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41396\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__41393\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__9009\ : Odrv12
    port map (
            O => \N__41390\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__41383\,
            I => \N__41380\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41374\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41374\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41374\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41365\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41365\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__41365\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__9001\ : CascadeMux
    port map (
            O => \N__41362\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__9000\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41356\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41356\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41347\
        );

    \I__8997\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41347\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__41347\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__41344\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__8994\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41338\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__41338\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__8990\ : Span4Mux_h
    port map (
            O => \N__41329\,
            I => \N__41325\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41328\,
            I => \N__41322\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__41325\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__41322\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__8986\ : CascadeMux
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41314\,
            I => \N__41311\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__41311\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41304\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__41307\,
            I => \N__41300\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__41304\,
            I => \N__41297\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41292\
        );

    \I__8979\ : InMux
    port map (
            O => \N__41300\,
            I => \N__41289\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__41297\,
            I => \N__41286\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41296\,
            I => \N__41281\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41295\,
            I => \N__41281\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__41292\,
            I => \N__41278\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41289\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__41286\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__41281\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__41278\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8970\ : IoInMux
    port map (
            O => \N__41269\,
            I => \N__41266\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41266\,
            I => \N__41263\
        );

    \I__8968\ : Span4Mux_s1_v
    port map (
            O => \N__41263\,
            I => \N__41234\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41223\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41223\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41260\,
            I => \N__41223\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41214\
        );

    \I__8963\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41214\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41214\
        );

    \I__8961\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41214\
        );

    \I__8960\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41205\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41254\,
            I => \N__41205\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41205\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41205\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41196\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41196\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41249\,
            I => \N__41196\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41196\
        );

    \I__8952\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41187\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41246\,
            I => \N__41187\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41187\
        );

    \I__8949\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41187\
        );

    \I__8948\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41178\
        );

    \I__8947\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41178\
        );

    \I__8946\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41178\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41240\,
            I => \N__41178\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41239\,
            I => \N__41171\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41238\,
            I => \N__41171\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41237\,
            I => \N__41171\
        );

    \I__8941\ : Span4Mux_v
    port map (
            O => \N__41234\,
            I => \N__41168\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41233\,
            I => \N__41159\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41159\
        );

    \I__8938\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41159\
        );

    \I__8937\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41159\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41156\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41145\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41145\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41196\,
            I => \N__41145\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41145\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__41178\,
            I => \N__41145\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41171\,
            I => \N__41142\
        );

    \I__8929\ : Sp12to4
    port map (
            O => \N__41168\,
            I => \N__41139\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__41159\,
            I => \N__41130\
        );

    \I__8927\ : Span4Mux_v
    port map (
            O => \N__41156\,
            I => \N__41130\
        );

    \I__8926\ : Span4Mux_v
    port map (
            O => \N__41145\,
            I => \N__41130\
        );

    \I__8925\ : Span4Mux_v
    port map (
            O => \N__41142\,
            I => \N__41130\
        );

    \I__8924\ : Span12Mux_h
    port map (
            O => \N__41139\,
            I => \N__41127\
        );

    \I__8923\ : Span4Mux_h
    port map (
            O => \N__41130\,
            I => \N__41124\
        );

    \I__8922\ : Span12Mux_v
    port map (
            O => \N__41127\,
            I => \N__41121\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__41124\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8920\ : Odrv12
    port map (
            O => \N__41121\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8919\ : InMux
    port map (
            O => \N__41116\,
            I => \N__41113\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41113\,
            I => \N__41110\
        );

    \I__8917\ : Sp12to4
    port map (
            O => \N__41110\,
            I => \N__41107\
        );

    \I__8916\ : Odrv12
    port map (
            O => \N__41107\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__8914\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41098\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__41098\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__41095\,
            I => \N__41092\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41092\,
            I => \N__41089\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41089\,
            I => \N__41086\
        );

    \I__8909\ : Odrv4
    port map (
            O => \N__41086\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__41083\,
            I => \N__41080\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41080\,
            I => \N__41077\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41077\,
            I => \N__41074\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__41074\,
            I => \N__41071\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__41071\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41062\
        );

    \I__8902\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41062\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__41062\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__41059\,
            I => \N__41055\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41050\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41050\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__41050\,
            I => \N__41046\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41043\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__41046\,
            I => \N__41040\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41043\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__41040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8892\ : CascadeMux
    port map (
            O => \N__41035\,
            I => \N__41032\
        );

    \I__8891\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41028\
        );

    \I__8890\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41025\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41019\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41019\
        );

    \I__8887\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41016\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__41019\,
            I => \N__41013\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__41016\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__41013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8883\ : InMux
    port map (
            O => \N__41008\,
            I => \N__41004\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41007\,
            I => \N__41001\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__41004\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__41001\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40993\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40990\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__40990\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40984\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40984\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__8874\ : CascadeMux
    port map (
            O => \N__40981\,
            I => \N__40978\
        );

    \I__8873\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40975\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40975\,
            I => \N__40972\
        );

    \I__8871\ : Odrv4
    port map (
            O => \N__40972\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40963\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40963\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40963\,
            I => \N__40959\
        );

    \I__8867\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40956\
        );

    \I__8866\ : Span4Mux_h
    port map (
            O => \N__40959\,
            I => \N__40953\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__40956\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__40953\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8863\ : CascadeMux
    port map (
            O => \N__40948\,
            I => \N__40945\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40939\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40944\,
            I => \N__40939\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40935\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40932\
        );

    \I__8858\ : Span4Mux_h
    port map (
            O => \N__40935\,
            I => \N__40929\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__40932\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__40929\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__40924\,
            I => \N__40921\
        );

    \I__8854\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40915\
        );

    \I__8853\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40915\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40915\,
            I => \N__40912\
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__40912\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40909\,
            I => \N__40906\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__40906\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__8848\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40900\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__40900\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40897\,
            I => \N__40894\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40894\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__8844\ : CascadeMux
    port map (
            O => \N__40891\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40885\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__40885\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40879\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40879\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__40876\,
            I => \N__40873\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40873\,
            I => \N__40870\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40870\,
            I => \N__40867\
        );

    \I__8836\ : Span4Mux_h
    port map (
            O => \N__40867\,
            I => \N__40864\
        );

    \I__8835\ : Odrv4
    port map (
            O => \N__40864\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__8834\ : CascadeMux
    port map (
            O => \N__40861\,
            I => \N__40857\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40852\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40852\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40852\,
            I => \N__40849\
        );

    \I__8830\ : Span4Mux_v
    port map (
            O => \N__40849\,
            I => \N__40845\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40842\
        );

    \I__8828\ : Span4Mux_v
    port map (
            O => \N__40845\,
            I => \N__40839\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__40842\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8826\ : Odrv4
    port map (
            O => \N__40839\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40834\,
            I => \N__40828\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40828\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40828\,
            I => \N__40824\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40827\,
            I => \N__40821\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__40824\,
            I => \N__40818\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__40821\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__40818\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8818\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__40810\,
            I => \N__40807\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__40807\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40804\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__8814\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40795\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40795\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__40795\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40792\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40789\,
            I => \N__40783\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40788\,
            I => \N__40779\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40774\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40774\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40771\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40768\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40763\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__40774\,
            I => \N__40763\
        );

    \I__8802\ : Span4Mux_v
    port map (
            O => \N__40771\,
            I => \N__40758\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__40768\,
            I => \N__40758\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__40763\,
            I => \N__40748\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__40758\,
            I => \N__40745\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__40757\,
            I => \N__40741\
        );

    \I__8797\ : CascadeMux
    port map (
            O => \N__40756\,
            I => \N__40737\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__40755\,
            I => \N__40733\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__40754\,
            I => \N__40729\
        );

    \I__8794\ : CascadeMux
    port map (
            O => \N__40753\,
            I => \N__40725\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__40752\,
            I => \N__40721\
        );

    \I__8792\ : CascadeMux
    port map (
            O => \N__40751\,
            I => \N__40717\
        );

    \I__8791\ : Span4Mux_h
    port map (
            O => \N__40748\,
            I => \N__40707\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__40745\,
            I => \N__40707\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40692\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40692\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40692\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40737\,
            I => \N__40692\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40692\
        );

    \I__8784\ : InMux
    port map (
            O => \N__40733\,
            I => \N__40692\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40692\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40675\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40675\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40725\,
            I => \N__40675\
        );

    \I__8779\ : InMux
    port map (
            O => \N__40724\,
            I => \N__40675\
        );

    \I__8778\ : InMux
    port map (
            O => \N__40721\,
            I => \N__40675\
        );

    \I__8777\ : InMux
    port map (
            O => \N__40720\,
            I => \N__40675\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40675\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40675\
        );

    \I__8774\ : CascadeMux
    port map (
            O => \N__40715\,
            I => \N__40672\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__40714\,
            I => \N__40668\
        );

    \I__8772\ : CascadeMux
    port map (
            O => \N__40713\,
            I => \N__40664\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__40712\,
            I => \N__40660\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__40707\,
            I => \N__40648\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40692\,
            I => \N__40648\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40648\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40672\,
            I => \N__40631\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40631\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40631\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40631\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40631\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40631\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40660\,
            I => \N__40631\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40631\
        );

    \I__8759\ : CascadeMux
    port map (
            O => \N__40658\,
            I => \N__40627\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__40657\,
            I => \N__40623\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__40656\,
            I => \N__40619\
        );

    \I__8756\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40613\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__40648\,
            I => \N__40600\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40631\,
            I => \N__40600\
        );

    \I__8753\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40585\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40585\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40585\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40585\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40585\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40585\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40585\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40580\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40580\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__40613\,
            I => \N__40566\
        );

    \I__8743\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40563\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40556\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40556\
        );

    \I__8740\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40556\
        );

    \I__8739\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40547\
        );

    \I__8738\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40547\
        );

    \I__8737\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40547\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40547\
        );

    \I__8735\ : Span4Mux_h
    port map (
            O => \N__40600\,
            I => \N__40539\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40585\,
            I => \N__40539\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40580\,
            I => \N__40539\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40534\
        );

    \I__8731\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40534\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40531\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40528\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40521\
        );

    \I__8727\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40521\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40521\
        );

    \I__8725\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40512\
        );

    \I__8724\ : InMux
    port map (
            O => \N__40571\,
            I => \N__40512\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40512\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40569\,
            I => \N__40512\
        );

    \I__8721\ : Span4Mux_v
    port map (
            O => \N__40566\,
            I => \N__40506\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__40563\,
            I => \N__40506\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__40556\,
            I => \N__40501\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__40547\,
            I => \N__40501\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40498\
        );

    \I__8716\ : Span4Mux_v
    port map (
            O => \N__40539\,
            I => \N__40494\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__40534\,
            I => \N__40489\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__40531\,
            I => \N__40489\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40528\,
            I => \N__40482\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40482\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40482\
        );

    \I__8710\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40479\
        );

    \I__8709\ : Span4Mux_v
    port map (
            O => \N__40506\,
            I => \N__40475\
        );

    \I__8708\ : Span4Mux_v
    port map (
            O => \N__40501\,
            I => \N__40470\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__40498\,
            I => \N__40470\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__40497\,
            I => \N__40466\
        );

    \I__8705\ : Span4Mux_v
    port map (
            O => \N__40494\,
            I => \N__40462\
        );

    \I__8704\ : Span12Mux_s11_h
    port map (
            O => \N__40489\,
            I => \N__40459\
        );

    \I__8703\ : Span4Mux_v
    port map (
            O => \N__40482\,
            I => \N__40456\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40479\,
            I => \N__40453\
        );

    \I__8701\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40450\
        );

    \I__8700\ : Span4Mux_s0_v
    port map (
            O => \N__40475\,
            I => \N__40445\
        );

    \I__8699\ : Span4Mux_v
    port map (
            O => \N__40470\,
            I => \N__40445\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40438\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40466\,
            I => \N__40438\
        );

    \I__8696\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40438\
        );

    \I__8695\ : Span4Mux_v
    port map (
            O => \N__40462\,
            I => \N__40435\
        );

    \I__8694\ : Span12Mux_v
    port map (
            O => \N__40459\,
            I => \N__40432\
        );

    \I__8693\ : Span4Mux_v
    port map (
            O => \N__40456\,
            I => \N__40427\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__40453\,
            I => \N__40427\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40450\,
            I => \N__40422\
        );

    \I__8690\ : Sp12to4
    port map (
            O => \N__40445\,
            I => \N__40422\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40419\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__40435\,
            I => \N__40416\
        );

    \I__8687\ : Span12Mux_v
    port map (
            O => \N__40432\,
            I => \N__40409\
        );

    \I__8686\ : Sp12to4
    port map (
            O => \N__40427\,
            I => \N__40409\
        );

    \I__8685\ : Span12Mux_s11_h
    port map (
            O => \N__40422\,
            I => \N__40409\
        );

    \I__8684\ : Span4Mux_v
    port map (
            O => \N__40419\,
            I => \N__40406\
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__40416\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8682\ : Odrv12
    port map (
            O => \N__40409\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__40406\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40399\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40396\,
            I => \N__40393\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40393\,
            I => \N__40390\
        );

    \I__8677\ : Odrv4
    port map (
            O => \N__40390\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40387\,
            I => \bfn_15_27_0_\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40379\
        );

    \I__8674\ : InMux
    port map (
            O => \N__40383\,
            I => \N__40376\
        );

    \I__8673\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40373\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__40379\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40376\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__40373\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8669\ : CascadeMux
    port map (
            O => \N__40366\,
            I => \N__40362\
        );

    \I__8668\ : InMux
    port map (
            O => \N__40365\,
            I => \N__40359\
        );

    \I__8667\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40356\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40359\,
            I => \N__40349\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__40356\,
            I => \N__40349\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40346\
        );

    \I__8663\ : InMux
    port map (
            O => \N__40354\,
            I => \N__40343\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__40349\,
            I => \N__40340\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40346\,
            I => \N__40337\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__40343\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__40340\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8658\ : Odrv12
    port map (
            O => \N__40337\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40330\,
            I => \N__40327\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__40327\,
            I => \N__40324\
        );

    \I__8655\ : Span4Mux_v
    port map (
            O => \N__40324\,
            I => \N__40321\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__40321\,
            I => \N__40318\
        );

    \I__8653\ : Sp12to4
    port map (
            O => \N__40318\,
            I => \N__40314\
        );

    \I__8652\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40311\
        );

    \I__8651\ : Odrv12
    port map (
            O => \N__40314\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40311\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40306\,
            I => \N__40303\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__40303\,
            I => \N__40300\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__8646\ : Sp12to4
    port map (
            O => \N__40297\,
            I => \N__40294\
        );

    \I__8645\ : Span12Mux_h
    port map (
            O => \N__40294\,
            I => \N__40291\
        );

    \I__8644\ : Odrv12
    port map (
            O => \N__40291\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__8643\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40285\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__8641\ : Span4Mux_v
    port map (
            O => \N__40282\,
            I => \N__40279\
        );

    \I__8640\ : Sp12to4
    port map (
            O => \N__40279\,
            I => \N__40276\
        );

    \I__8639\ : Odrv12
    port map (
            O => \N__40276\,
            I => \pwm_generator_inst.O_12\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40273\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__8637\ : InMux
    port map (
            O => \N__40270\,
            I => \N__40267\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__40267\,
            I => \N__40264\
        );

    \I__8635\ : Sp12to4
    port map (
            O => \N__40264\,
            I => \N__40261\
        );

    \I__8634\ : Span12Mux_s6_v
    port map (
            O => \N__40261\,
            I => \N__40258\
        );

    \I__8633\ : Odrv12
    port map (
            O => \N__40258\,
            I => \pwm_generator_inst.O_13\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40255\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40252\,
            I => \N__40249\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__40249\,
            I => \N__40246\
        );

    \I__8629\ : Span12Mux_s6_v
    port map (
            O => \N__40246\,
            I => \N__40243\
        );

    \I__8628\ : Odrv12
    port map (
            O => \N__40243\,
            I => \pwm_generator_inst.O_14\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40240\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40237\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40234\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__40231\,
            I => \N__40228\
        );

    \I__8623\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40224\
        );

    \I__8622\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40221\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__40224\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__40221\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40213\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40209\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40206\
        );

    \I__8616\ : Odrv4
    port map (
            O => \N__40209\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40206\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__40201\,
            I => \N__40197\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40194\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40191\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__40194\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40191\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40186\,
            I => \N__40183\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__40183\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40174\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40179\,
            I => \N__40174\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40174\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40168\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40168\,
            I => \N__40164\
        );

    \I__8602\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40161\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40164\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__40161\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__40156\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40153\,
            I => \N__40150\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40150\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__40147\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__8595\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40141\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40141\,
            I => \N__40138\
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__40138\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40126\
        );

    \I__8590\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40126\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40126\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40123\,
            I => \N__40120\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40120\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40114\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40114\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__8584\ : CascadeMux
    port map (
            O => \N__40111\,
            I => \N__40108\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40108\,
            I => \N__40102\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40102\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40102\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__40099\,
            I => \N__40095\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40090\
        );

    \I__8578\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40090\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__40090\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40087\,
            I => \N__40084\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40084\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40075\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40075\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__40075\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__8571\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40068\
        );

    \I__8570\ : InMux
    port map (
            O => \N__40071\,
            I => \N__40065\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__40068\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__40065\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__8567\ : CascadeMux
    port map (
            O => \N__40060\,
            I => \N__40057\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40051\
        );

    \I__8565\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40051\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40051\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40048\,
            I => \N__40044\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40047\,
            I => \N__40041\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__40044\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__40041\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__40036\,
            I => \N__40032\
        );

    \I__8558\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40028\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40032\,
            I => \N__40023\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40031\,
            I => \N__40023\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__40028\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__40023\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__40018\,
            I => \N__40015\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40015\,
            I => \N__40010\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40014\,
            I => \N__40005\
        );

    \I__8550\ : InMux
    port map (
            O => \N__40013\,
            I => \N__40005\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__40010\,
            I => \N__40000\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__40005\,
            I => \N__40000\
        );

    \I__8547\ : Span4Mux_h
    port map (
            O => \N__40000\,
            I => \N__39997\
        );

    \I__8546\ : Span4Mux_v
    port map (
            O => \N__39997\,
            I => \N__39993\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39990\
        );

    \I__8544\ : Span4Mux_v
    port map (
            O => \N__39993\,
            I => \N__39987\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__39990\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__39987\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39978\
        );

    \I__8540\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39975\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__39978\,
            I => \N__39972\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39975\,
            I => \N__39969\
        );

    \I__8537\ : Span4Mux_h
    port map (
            O => \N__39972\,
            I => \N__39966\
        );

    \I__8536\ : Span4Mux_s3_h
    port map (
            O => \N__39969\,
            I => \N__39963\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__39966\,
            I => \N__39960\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__39963\,
            I => \N__39957\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__39960\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__39957\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39952\,
            I => \N__39949\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__39949\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__39946\,
            I => \N__39943\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39943\,
            I => \N__39939\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__39942\,
            I => \N__39936\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__39939\,
            I => \N__39933\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39929\
        );

    \I__8524\ : Span4Mux_v
    port map (
            O => \N__39933\,
            I => \N__39926\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39923\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39920\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__39926\,
            I => \N__39917\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__39923\,
            I => \N__39912\
        );

    \I__8519\ : Span4Mux_v
    port map (
            O => \N__39920\,
            I => \N__39907\
        );

    \I__8518\ : Span4Mux_h
    port map (
            O => \N__39917\,
            I => \N__39907\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39916\,
            I => \N__39904\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39901\
        );

    \I__8515\ : Span12Mux_v
    port map (
            O => \N__39912\,
            I => \N__39898\
        );

    \I__8514\ : Span4Mux_v
    port map (
            O => \N__39907\,
            I => \N__39893\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39904\,
            I => \N__39893\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8511\ : Odrv12
    port map (
            O => \N__39898\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8510\ : Odrv4
    port map (
            O => \N__39893\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__39886\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39877\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39882\,
            I => \N__39877\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__39877\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39868\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39868\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39868\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39865\,
            I => \N__39859\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39859\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39859\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__8499\ : CascadeMux
    port map (
            O => \N__39856\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39847\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39852\,
            I => \N__39847\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__39847\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__39844\,
            I => \N__39841\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39837\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39834\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__39837\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39834\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39829\,
            I => \N__39823\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39823\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39823\,
            I => \N__39819\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39816\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__39819\,
            I => \N__39813\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39816\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__8484\ : Odrv4
    port map (
            O => \N__39813\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39808\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__39805\,
            I => \N__39801\
        );

    \I__8481\ : CascadeMux
    port map (
            O => \N__39804\,
            I => \N__39798\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39793\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39793\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39789\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39786\
        );

    \I__8476\ : Span4Mux_h
    port map (
            O => \N__39789\,
            I => \N__39783\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39786\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__39783\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39778\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__39775\,
            I => \N__39772\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39766\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39771\,
            I => \N__39766\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39766\,
            I => \N__39762\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39759\
        );

    \I__8467\ : Span4Mux_h
    port map (
            O => \N__39762\,
            I => \N__39756\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39759\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__39756\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39751\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39742\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39747\,
            I => \N__39742\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39742\,
            I => \N__39738\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39741\,
            I => \N__39735\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__39738\,
            I => \N__39732\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__39735\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__39732\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39727\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__39724\,
            I => \N__39720\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39723\,
            I => \N__39717\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39714\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39717\,
            I => \N__39708\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39714\,
            I => \N__39708\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39713\,
            I => \N__39705\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__39708\,
            I => \N__39702\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39705\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__39702\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39697\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39694\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__39691\,
            I => \N__39688\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39688\,
            I => \N__39684\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39681\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39677\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39681\,
            I => \N__39674\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39671\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__39677\,
            I => \N__39668\
        );

    \I__8437\ : Span12Mux_v
    port map (
            O => \N__39674\,
            I => \N__39665\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39671\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8435\ : Odrv4
    port map (
            O => \N__39668\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8434\ : Odrv12
    port map (
            O => \N__39665\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39655\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39655\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39652\,
            I => \bfn_15_14_0_\
        );

    \I__8430\ : InMux
    port map (
            O => \N__39649\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39646\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__8428\ : InMux
    port map (
            O => \N__39643\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39640\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39631\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39636\,
            I => \N__39631\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39631\,
            I => \N__39627\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39630\,
            I => \N__39624\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__39627\,
            I => \N__39621\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__39624\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__39621\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39616\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__39613\,
            I => \N__39609\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39604\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39604\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39604\,
            I => \N__39600\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39603\,
            I => \N__39597\
        );

    \I__8413\ : Span12Mux_s7_v
    port map (
            O => \N__39600\,
            I => \N__39594\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39597\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8411\ : Odrv12
    port map (
            O => \N__39594\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39589\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39581\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39576\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39584\,
            I => \N__39576\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39581\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39576\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__8404\ : InMux
    port map (
            O => \N__39571\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39561\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39561\
        );

    \I__8401\ : InMux
    port map (
            O => \N__39566\,
            I => \N__39558\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__39561\,
            I => \N__39555\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39558\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__39555\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39550\,
            I => \bfn_15_15_0_\
        );

    \I__8396\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39543\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39540\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39537\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__39540\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8392\ : Odrv4
    port map (
            O => \N__39537\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39532\,
            I => \bfn_15_13_0_\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39525\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39528\,
            I => \N__39522\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__39525\,
            I => \N__39519\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39522\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__39519\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39514\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__8384\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39507\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39504\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__39507\,
            I => \N__39501\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__39504\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8380\ : Odrv4
    port map (
            O => \N__39501\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39496\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39493\,
            I => \N__39489\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39486\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__39489\,
            I => \N__39483\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39486\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8374\ : Odrv4
    port map (
            O => \N__39483\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39478\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39471\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39474\,
            I => \N__39468\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__39471\,
            I => \N__39465\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39468\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8368\ : Odrv4
    port map (
            O => \N__39465\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39460\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39454\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__39454\,
            I => \N__39450\
        );

    \I__8364\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39447\
        );

    \I__8363\ : Span4Mux_v
    port map (
            O => \N__39450\,
            I => \N__39444\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__39447\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__39444\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39439\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39432\
        );

    \I__8358\ : InMux
    port map (
            O => \N__39435\,
            I => \N__39429\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__39432\,
            I => \N__39426\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39429\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8355\ : Odrv12
    port map (
            O => \N__39426\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8354\ : InMux
    port map (
            O => \N__39421\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39418\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39415\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__39412\,
            I => \N__39409\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39409\,
            I => \N__39404\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39408\,
            I => \N__39401\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__39407\,
            I => \N__39398\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__39404\,
            I => \N__39393\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39401\,
            I => \N__39393\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39390\
        );

    \I__8344\ : Span4Mux_v
    port map (
            O => \N__39393\,
            I => \N__39387\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39390\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__39387\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39378\
        );

    \I__8340\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39375\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39372\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__39375\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8337\ : Odrv12
    port map (
            O => \N__39372\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8336\ : InMux
    port map (
            O => \N__39367\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39360\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39357\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39360\,
            I => \N__39354\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__39357\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__39354\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39349\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39346\,
            I => \N__39342\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39345\,
            I => \N__39339\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__39342\,
            I => \N__39336\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__39339\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8325\ : Odrv4
    port map (
            O => \N__39336\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39331\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39324\
        );

    \I__8322\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39321\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__39324\,
            I => \N__39318\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__39321\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8319\ : Odrv4
    port map (
            O => \N__39318\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8318\ : InMux
    port map (
            O => \N__39313\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__8317\ : InMux
    port map (
            O => \N__39310\,
            I => \N__39306\
        );

    \I__8316\ : InMux
    port map (
            O => \N__39309\,
            I => \N__39303\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39306\,
            I => \N__39300\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__39303\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__39300\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39295\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__8311\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39288\
        );

    \I__8310\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39285\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__39288\,
            I => \N__39282\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__39285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8307\ : Odrv12
    port map (
            O => \N__39282\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39277\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__8305\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39270\
        );

    \I__8304\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39267\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39264\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39267\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8301\ : Odrv12
    port map (
            O => \N__39264\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39259\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39256\,
            I => \N__39253\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39253\,
            I => \N__39250\
        );

    \I__8297\ : Odrv12
    port map (
            O => \N__39250\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__39247\,
            I => \N__39244\
        );

    \I__8295\ : InMux
    port map (
            O => \N__39244\,
            I => \N__39241\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__8293\ : Span4Mux_v
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__8292\ : Odrv4
    port map (
            O => \N__39235\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__8291\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39229\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__39229\,
            I => \N__39226\
        );

    \I__8289\ : Odrv4
    port map (
            O => \N__39226\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__8288\ : CascadeMux
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__8287\ : InMux
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__39217\,
            I => \N__39214\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__39214\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__8284\ : InMux
    port map (
            O => \N__39211\,
            I => \N__39208\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__39208\,
            I => \N__39205\
        );

    \I__8282\ : Odrv12
    port map (
            O => \N__39205\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__39202\,
            I => \N__39199\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39196\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39196\,
            I => \N__39193\
        );

    \I__8278\ : Odrv12
    port map (
            O => \N__39193\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__8277\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39187\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39187\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__39184\,
            I => \N__39181\
        );

    \I__8274\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39178\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__39178\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39172\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39172\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__8270\ : CascadeMux
    port map (
            O => \N__39169\,
            I => \N__39166\
        );

    \I__8269\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39163\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__39160\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39154\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__39154\,
            I => \N__39151\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__39151\,
            I => \N__39148\
        );

    \I__8263\ : Odrv4
    port map (
            O => \N__39148\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__39145\,
            I => \N__39142\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39139\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__39139\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8259\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39133\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__39133\,
            I => \N__39130\
        );

    \I__8257\ : Odrv12
    port map (
            O => \N__39130\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39121\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__39121\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__39118\,
            I => \N__39115\
        );

    \I__8252\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39112\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__39112\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8250\ : CascadeMux
    port map (
            O => \N__39109\,
            I => \N__39106\
        );

    \I__8249\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39103\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39103\,
            I => \N__39100\
        );

    \I__8247\ : Odrv12
    port map (
            O => \N__39100\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39094\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__39094\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8244\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39088\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__39088\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__39085\,
            I => \N__39082\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39079\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39076\
        );

    \I__8239\ : Odrv4
    port map (
            O => \N__39076\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__8238\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39070\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__39070\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__39067\,
            I => \N__39064\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39061\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__39061\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8233\ : InMux
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__39055\,
            I => \N__39052\
        );

    \I__8231\ : Odrv12
    port map (
            O => \N__39052\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__39049\,
            I => \N__39046\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39043\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__39043\,
            I => \N__39040\
        );

    \I__8227\ : Odrv4
    port map (
            O => \N__39040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8226\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39034\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__39031\,
            I => \N__39028\
        );

    \I__8223\ : InMux
    port map (
            O => \N__39028\,
            I => \N__39025\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__39025\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__39022\,
            I => \N__39019\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39016\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__39016\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__8218\ : InMux
    port map (
            O => \N__39013\,
            I => \N__39010\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__39010\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8216\ : InMux
    port map (
            O => \N__39007\,
            I => \N__39004\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__39004\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__39001\,
            I => \N__38998\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38998\,
            I => \N__38995\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38992\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__38992\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8210\ : InMux
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38986\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__38983\,
            I => \N__38980\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38977\,
            I => \N__38974\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__38974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38968\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38959\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38953\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__38953\,
            I => \N__38950\
        );

    \I__8197\ : Odrv12
    port map (
            O => \N__38950\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__38947\,
            I => \N__38944\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38941\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38941\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38932\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38932\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38932\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__38929\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38923\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38923\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__8187\ : IoInMux
    port map (
            O => \N__38920\,
            I => \N__38917\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38917\,
            I => \N__38914\
        );

    \I__8185\ : Span4Mux_s2_v
    port map (
            O => \N__38914\,
            I => \N__38911\
        );

    \I__8184\ : Span4Mux_h
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__38908\,
            I => s4_phy_c
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__38905\,
            I => \N__38902\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38896\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__38896\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38893\,
            I => \N__38890\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38890\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__8176\ : InMux
    port map (
            O => \N__38887\,
            I => \N__38884\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__38884\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__38881\,
            I => \N__38878\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38875\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38875\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__38872\,
            I => \N__38869\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38866\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__38866\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38863\,
            I => \N__38860\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38860\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__8166\ : CascadeMux
    port map (
            O => \N__38857\,
            I => \N__38854\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38854\,
            I => \N__38851\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38851\,
            I => \N__38848\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38848\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38842\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38842\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__38839\,
            I => \N__38836\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38833\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38833\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38827\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38827\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38821\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38821\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__8153\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38815\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__38815\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38809\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__38809\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38806\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38803\,
            I => \N__38794\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38794\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38787\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38774\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38799\,
            I => \N__38771\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__38794\,
            I => \N__38768\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38759\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38759\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38791\,
            I => \N__38759\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38759\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38787\,
            I => \N__38756\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38745\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38785\,
            I => \N__38745\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38745\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38745\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38745\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38781\,
            I => \N__38742\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38739\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38721\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38778\,
            I => \N__38721\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38721\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38774\,
            I => \N__38712\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38771\,
            I => \N__38712\
        );

    \I__8125\ : Span4Mux_h
    port map (
            O => \N__38768\,
            I => \N__38712\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38759\,
            I => \N__38712\
        );

    \I__8123\ : Sp12to4
    port map (
            O => \N__38756\,
            I => \N__38709\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__38745\,
            I => \N__38703\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38703\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38739\,
            I => \N__38700\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38694\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38694\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38683\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38683\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38683\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38683\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38683\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38731\,
            I => \N__38674\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38674\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38674\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38728\,
            I => \N__38674\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__38721\,
            I => \N__38671\
        );

    \I__8107\ : Span4Mux_v
    port map (
            O => \N__38712\,
            I => \N__38668\
        );

    \I__8106\ : Span12Mux_h
    port map (
            O => \N__38709\,
            I => \N__38665\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38662\
        );

    \I__8104\ : Span4Mux_h
    port map (
            O => \N__38703\,
            I => \N__38657\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__38700\,
            I => \N__38657\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38654\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__38694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38683\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38674\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8098\ : Odrv4
    port map (
            O => \N__38671\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__38668\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8096\ : Odrv12
    port map (
            O => \N__38665\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__38662\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__38657\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38654\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38635\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38632\,
            I => \N__38629\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38629\,
            I => \N__38626\
        );

    \I__8089\ : Span4Mux_h
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__8088\ : Span4Mux_h
    port map (
            O => \N__38623\,
            I => \N__38620\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__38620\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38614\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38614\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38608\,
            I => \N__38605\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__38605\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__38602\,
            I => \N__38599\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38596\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__38596\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38590\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38590\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__38584\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__38581\,
            I => \N__38578\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38575\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__38575\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__38572\,
            I => \N__38569\
        );

    \I__8070\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38566\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38560\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__38560\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38554\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__38554\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__38551\,
            I => \N__38548\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38545\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__38542\,
            I => \N__38539\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38539\,
            I => \N__38536\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38536\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__8056\ : Span4Mux_v
    port map (
            O => \N__38527\,
            I => \N__38524\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__38524\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38515\,
            I => \N__38512\
        );

    \I__8051\ : Span4Mux_v
    port map (
            O => \N__38512\,
            I => \N__38508\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38505\
        );

    \I__8049\ : Span4Mux_v
    port map (
            O => \N__38508\,
            I => \N__38500\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38497\
        );

    \I__8047\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38494\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38491\
        );

    \I__8045\ : Sp12to4
    port map (
            O => \N__38500\,
            I => \N__38488\
        );

    \I__8044\ : Span4Mux_v
    port map (
            O => \N__38497\,
            I => \N__38485\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38494\,
            I => \N__38482\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__38491\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8041\ : Odrv12
    port map (
            O => \N__38488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__38485\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8039\ : Odrv4
    port map (
            O => \N__38482\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38473\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38467\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__38467\,
            I => \N__38464\
        );

    \I__8035\ : Odrv4
    port map (
            O => \N__38464\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__38461\,
            I => \N__38458\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38455\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__38455\,
            I => \N__38452\
        );

    \I__8031\ : Span4Mux_h
    port map (
            O => \N__38452\,
            I => \N__38449\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__38449\,
            I => \N__38444\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38441\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__38447\,
            I => \N__38438\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__38444\,
            I => \N__38434\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__38441\,
            I => \N__38431\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38438\,
            I => \N__38428\
        );

    \I__8024\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38425\
        );

    \I__8023\ : Span4Mux_v
    port map (
            O => \N__38434\,
            I => \N__38422\
        );

    \I__8022\ : Span4Mux_v
    port map (
            O => \N__38431\,
            I => \N__38417\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38428\,
            I => \N__38417\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__38425\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__38422\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__38417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38410\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__8016\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38404\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38404\,
            I => \N__38401\
        );

    \I__8014\ : Odrv12
    port map (
            O => \N__38401\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__8013\ : CascadeMux
    port map (
            O => \N__38398\,
            I => \N__38395\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38389\
        );

    \I__8010\ : Sp12to4
    port map (
            O => \N__38389\,
            I => \N__38385\
        );

    \I__8009\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38380\
        );

    \I__8008\ : Span12Mux_v
    port map (
            O => \N__38385\,
            I => \N__38377\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38384\,
            I => \N__38374\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38383\,
            I => \N__38371\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__38380\,
            I => \N__38368\
        );

    \I__8004\ : Odrv12
    port map (
            O => \N__38377\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38374\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38371\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__38368\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__8000\ : InMux
    port map (
            O => \N__38359\,
            I => \bfn_14_20_0_\
        );

    \I__7999\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38353\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__38353\,
            I => \N__38350\
        );

    \I__7997\ : Odrv12
    port map (
            O => \N__38350\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__38347\,
            I => \N__38344\
        );

    \I__7995\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38341\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38341\,
            I => \N__38338\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__38338\,
            I => \N__38334\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38330\
        );

    \I__7991\ : Sp12to4
    port map (
            O => \N__38334\,
            I => \N__38326\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38333\,
            I => \N__38323\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38330\,
            I => \N__38320\
        );

    \I__7988\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38317\
        );

    \I__7987\ : Span12Mux_h
    port map (
            O => \N__38326\,
            I => \N__38314\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38323\,
            I => \N__38311\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__38320\,
            I => \N__38308\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__38317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7983\ : Odrv12
    port map (
            O => \N__38314\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__38311\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__38308\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__7980\ : InMux
    port map (
            O => \N__38299\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38293\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38293\,
            I => \N__38290\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__38290\,
            I => \N__38287\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__38287\,
            I => \N__38284\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__38284\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__7974\ : CascadeMux
    port map (
            O => \N__38281\,
            I => \N__38278\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__7971\ : Span4Mux_v
    port map (
            O => \N__38272\,
            I => \N__38268\
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__38271\,
            I => \N__38265\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__38268\,
            I => \N__38261\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38258\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__38264\,
            I => \N__38254\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__38261\,
            I => \N__38249\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__38258\,
            I => \N__38249\
        );

    \I__7964\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38246\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38243\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__38249\,
            I => \N__38240\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__38246\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__38243\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__38240\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38233\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38224\
        );

    \I__7955\ : Span4Mux_v
    port map (
            O => \N__38224\,
            I => \N__38221\
        );

    \I__7954\ : Span4Mux_h
    port map (
            O => \N__38221\,
            I => \N__38217\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38220\,
            I => \N__38214\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__38217\,
            I => \N__38207\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__38214\,
            I => \N__38207\
        );

    \I__7950\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38204\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38201\
        );

    \I__7948\ : Span4Mux_h
    port map (
            O => \N__38207\,
            I => \N__38198\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__38204\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__38201\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__38198\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__38191\,
            I => \N__38188\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__38185\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38182\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38176\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38176\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__38173\,
            I => \N__38170\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38167\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__7935\ : Span4Mux_v
    port map (
            O => \N__38164\,
            I => \N__38161\
        );

    \I__7934\ : Span4Mux_h
    port map (
            O => \N__38161\,
            I => \N__38158\
        );

    \I__7933\ : Span4Mux_h
    port map (
            O => \N__38158\,
            I => \N__38153\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38149\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38146\
        );

    \I__7930\ : Span4Mux_h
    port map (
            O => \N__38153\,
            I => \N__38143\
        );

    \I__7929\ : InMux
    port map (
            O => \N__38152\,
            I => \N__38140\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__38149\,
            I => \N__38137\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38146\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__38143\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__38140\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__38137\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__7923\ : InMux
    port map (
            O => \N__38128\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__7922\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__7919\ : Span4Mux_h
    port map (
            O => \N__38116\,
            I => \N__38113\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__38113\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__7917\ : CascadeMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__7916\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38101\
        );

    \I__7914\ : Span4Mux_v
    port map (
            O => \N__38101\,
            I => \N__38097\
        );

    \I__7913\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38094\
        );

    \I__7912\ : Sp12to4
    port map (
            O => \N__38097\,
            I => \N__38089\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__38094\,
            I => \N__38086\
        );

    \I__7910\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38083\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38080\
        );

    \I__7908\ : Span12Mux_h
    port map (
            O => \N__38089\,
            I => \N__38077\
        );

    \I__7907\ : Span4Mux_v
    port map (
            O => \N__38086\,
            I => \N__38074\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__38071\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__38080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7904\ : Odrv12
    port map (
            O => \N__38077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7903\ : Odrv4
    port map (
            O => \N__38074\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__38071\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38062\,
            I => \N__38059\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38059\,
            I => \N__38056\
        );

    \I__7899\ : Span4Mux_h
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__7898\ : Span4Mux_h
    port map (
            O => \N__38053\,
            I => \N__38050\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__38050\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__7896\ : CascadeMux
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38041\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__38041\,
            I => \N__38037\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38040\,
            I => \N__38033\
        );

    \I__7892\ : Span4Mux_h
    port map (
            O => \N__38037\,
            I => \N__38030\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38026\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__38033\,
            I => \N__38023\
        );

    \I__7889\ : Sp12to4
    port map (
            O => \N__38030\,
            I => \N__38020\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38017\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38014\
        );

    \I__7886\ : Span4Mux_v
    port map (
            O => \N__38023\,
            I => \N__38011\
        );

    \I__7885\ : Span12Mux_v
    port map (
            O => \N__38020\,
            I => \N__38006\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__38017\,
            I => \N__38006\
        );

    \I__7883\ : Odrv12
    port map (
            O => \N__38014\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__38011\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7881\ : Odrv12
    port map (
            O => \N__38006\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37999\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37993\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37993\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__37990\,
            I => \N__37987\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37987\,
            I => \N__37984\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37984\,
            I => \N__37980\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__37983\,
            I => \N__37977\
        );

    \I__7873\ : Span4Mux_v
    port map (
            O => \N__37980\,
            I => \N__37972\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37977\,
            I => \N__37969\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37966\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37963\
        );

    \I__7869\ : Span4Mux_h
    port map (
            O => \N__37972\,
            I => \N__37960\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37957\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37952\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37952\
        );

    \I__7865\ : Span4Mux_h
    port map (
            O => \N__37960\,
            I => \N__37947\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__37957\,
            I => \N__37947\
        );

    \I__7863\ : Odrv12
    port map (
            O => \N__37952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__37947\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7861\ : InMux
    port map (
            O => \N__37942\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__7860\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37936\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__37936\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__37933\,
            I => \N__37930\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37930\,
            I => \N__37927\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37927\,
            I => \N__37921\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__37926\,
            I => \N__37918\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37915\
        );

    \I__7853\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37912\
        );

    \I__7852\ : Span12Mux_v
    port map (
            O => \N__37921\,
            I => \N__37909\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37906\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37915\,
            I => \N__37903\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37900\
        );

    \I__7848\ : Odrv12
    port map (
            O => \N__37909\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__37906\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7846\ : Odrv12
    port map (
            O => \N__37903\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__37900\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37891\,
            I => \bfn_14_19_0_\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37885\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37882\
        );

    \I__7841\ : Sp12to4
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__7840\ : Span12Mux_v
    port map (
            O => \N__37879\,
            I => \N__37873\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37870\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37867\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37864\
        );

    \I__7836\ : Span12Mux_h
    port map (
            O => \N__37873\,
            I => \N__37859\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37859\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37856\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37864\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__7832\ : Odrv12
    port map (
            O => \N__37859\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__37856\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37843\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37843\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37840\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37834\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37834\,
            I => \N__37831\
        );

    \I__7824\ : Sp12to4
    port map (
            O => \N__37831\,
            I => \N__37827\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37824\
        );

    \I__7822\ : Span12Mux_v
    port map (
            O => \N__37827\,
            I => \N__37819\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37824\,
            I => \N__37816\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37813\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37810\
        );

    \I__7818\ : Span12Mux_h
    port map (
            O => \N__37819\,
            I => \N__37807\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__37816\,
            I => \N__37802\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37802\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__37810\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7814\ : Odrv12
    port map (
            O => \N__37807\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__37802\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7812\ : CascadeMux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37789\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37789\,
            I => \N__37786\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__37786\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37783\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37777\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37777\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__37774\,
            I => \N__37771\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37768\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__37768\,
            I => \N__37765\
        );

    \I__7802\ : Span4Mux_v
    port map (
            O => \N__37765\,
            I => \N__37759\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37756\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37753\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37750\
        );

    \I__7798\ : Sp12to4
    port map (
            O => \N__37759\,
            I => \N__37747\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37756\,
            I => \N__37742\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__37753\,
            I => \N__37742\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37739\
        );

    \I__7794\ : Span12Mux_h
    port map (
            O => \N__37747\,
            I => \N__37736\
        );

    \I__7793\ : Span4Mux_v
    port map (
            O => \N__37742\,
            I => \N__37733\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__37739\,
            I => \N__37730\
        );

    \I__7791\ : Odrv12
    port map (
            O => \N__37736\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__37733\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7789\ : Odrv4
    port map (
            O => \N__37730\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37723\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37717\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37714\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__37714\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__7784\ : CascadeMux
    port map (
            O => \N__37711\,
            I => \N__37708\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37705\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37700\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37696\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37693\
        );

    \I__7779\ : Span12Mux_v
    port map (
            O => \N__37700\,
            I => \N__37690\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37699\,
            I => \N__37687\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37696\,
            I => \N__37682\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37682\
        );

    \I__7775\ : Odrv12
    port map (
            O => \N__37690\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37687\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__37682\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37675\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37672\,
            I => \N__37669\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37669\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__7769\ : CascadeMux
    port map (
            O => \N__37666\,
            I => \N__37663\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37663\,
            I => \N__37660\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__37660\,
            I => \N__37657\
        );

    \I__7766\ : Sp12to4
    port map (
            O => \N__37657\,
            I => \N__37652\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__37656\,
            I => \N__37649\
        );

    \I__7764\ : CascadeMux
    port map (
            O => \N__37655\,
            I => \N__37646\
        );

    \I__7763\ : Span12Mux_v
    port map (
            O => \N__37652\,
            I => \N__37642\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37639\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37636\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37645\,
            I => \N__37633\
        );

    \I__7759\ : Span12Mux_h
    port map (
            O => \N__37642\,
            I => \N__37628\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37639\,
            I => \N__37628\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37636\,
            I => \N__37625\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37633\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__37628\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__37625\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37618\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37612\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37612\,
            I => \N__37609\
        );

    \I__7750\ : Odrv12
    port map (
            O => \N__37609\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__37606\,
            I => \N__37603\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37600\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37597\
        );

    \I__7746\ : Span4Mux_h
    port map (
            O => \N__37597\,
            I => \N__37594\
        );

    \I__7745\ : Span4Mux_h
    port map (
            O => \N__37594\,
            I => \N__37589\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37593\,
            I => \N__37586\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37592\,
            I => \N__37583\
        );

    \I__7742\ : Span4Mux_v
    port map (
            O => \N__37589\,
            I => \N__37577\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__37586\,
            I => \N__37577\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__37583\,
            I => \N__37574\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37571\
        );

    \I__7738\ : Span4Mux_h
    port map (
            O => \N__37577\,
            I => \N__37568\
        );

    \I__7737\ : Span4Mux_v
    port map (
            O => \N__37574\,
            I => \N__37565\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37571\,
            I => \N__37560\
        );

    \I__7735\ : Span4Mux_v
    port map (
            O => \N__37568\,
            I => \N__37560\
        );

    \I__7734\ : Odrv4
    port map (
            O => \N__37565\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__37560\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37555\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__7731\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37549\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__37549\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__37546\,
            I => \N__37543\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37543\,
            I => \N__37540\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__37540\,
            I => \N__37537\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__37537\,
            I => \N__37531\
        );

    \I__7725\ : InMux
    port map (
            O => \N__37536\,
            I => \N__37528\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37525\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37522\
        );

    \I__7722\ : Sp12to4
    port map (
            O => \N__37531\,
            I => \N__37519\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__37528\,
            I => \N__37514\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__37525\,
            I => \N__37514\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37522\,
            I => \N__37511\
        );

    \I__7718\ : Span12Mux_v
    port map (
            O => \N__37519\,
            I => \N__37508\
        );

    \I__7717\ : Span4Mux_v
    port map (
            O => \N__37514\,
            I => \N__37503\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__37511\,
            I => \N__37503\
        );

    \I__7715\ : Odrv12
    port map (
            O => \N__37508\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__7714\ : Odrv4
    port map (
            O => \N__37503\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37498\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37492\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__37492\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__37489\,
            I => \N__37486\
        );

    \I__7709\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37483\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37483\,
            I => \N__37479\
        );

    \I__7707\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37476\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__37479\,
            I => \N__37472\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37468\
        );

    \I__7704\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37465\
        );

    \I__7703\ : Span4Mux_v
    port map (
            O => \N__37472\,
            I => \N__37462\
        );

    \I__7702\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37459\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__37468\,
            I => \N__37456\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__37465\,
            I => \N__37453\
        );

    \I__7699\ : Sp12to4
    port map (
            O => \N__37462\,
            I => \N__37450\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37459\,
            I => \N__37447\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__37456\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7696\ : Odrv12
    port map (
            O => \N__37453\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7695\ : Odrv12
    port map (
            O => \N__37450\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7694\ : Odrv4
    port map (
            O => \N__37447\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7693\ : InMux
    port map (
            O => \N__37438\,
            I => \bfn_14_18_0_\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37431\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__37434\,
            I => \N__37428\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37424\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37421\
        );

    \I__7688\ : CascadeMux
    port map (
            O => \N__37427\,
            I => \N__37418\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__37424\,
            I => \N__37415\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__37421\,
            I => \N__37411\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37408\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__37415\,
            I => \N__37405\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37414\,
            I => \N__37402\
        );

    \I__7682\ : Span4Mux_h
    port map (
            O => \N__37411\,
            I => \N__37397\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37408\,
            I => \N__37397\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__37405\,
            I => \N__37394\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37402\,
            I => \N__37391\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__37397\,
            I => \N__37388\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__37394\,
            I => \N__37383\
        );

    \I__7676\ : Span4Mux_v
    port map (
            O => \N__37391\,
            I => \N__37383\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__37388\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__37383\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__7673\ : CascadeMux
    port map (
            O => \N__37378\,
            I => \N__37375\
        );

    \I__7672\ : InMux
    port map (
            O => \N__37375\,
            I => \N__37372\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__37372\,
            I => \N__37369\
        );

    \I__7670\ : Odrv12
    port map (
            O => \N__37369\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37366\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__7668\ : InMux
    port map (
            O => \N__37363\,
            I => \N__37360\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__37360\,
            I => \N__37357\
        );

    \I__7666\ : Span4Mux_h
    port map (
            O => \N__37357\,
            I => \N__37354\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__37354\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__7664\ : CascadeMux
    port map (
            O => \N__37351\,
            I => \N__37348\
        );

    \I__7663\ : InMux
    port map (
            O => \N__37348\,
            I => \N__37345\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__37345\,
            I => \N__37342\
        );

    \I__7661\ : Span4Mux_v
    port map (
            O => \N__37342\,
            I => \N__37337\
        );

    \I__7660\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37334\
        );

    \I__7659\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37331\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__37337\,
            I => \N__37327\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37324\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37321\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37318\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__37327\,
            I => \N__37313\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__37324\,
            I => \N__37313\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__37321\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__37318\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__37313\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37306\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__37300\,
            I => \N__37297\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__37297\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__7645\ : CascadeMux
    port map (
            O => \N__37294\,
            I => \N__37291\
        );

    \I__7644\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37288\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37288\,
            I => \N__37284\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37280\
        );

    \I__7641\ : Span4Mux_v
    port map (
            O => \N__37284\,
            I => \N__37277\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37274\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37271\
        );

    \I__7638\ : Span4Mux_h
    port map (
            O => \N__37277\,
            I => \N__37268\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37264\
        );

    \I__7636\ : Span4Mux_h
    port map (
            O => \N__37271\,
            I => \N__37259\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__37268\,
            I => \N__37259\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37267\,
            I => \N__37256\
        );

    \I__7633\ : Span4Mux_v
    port map (
            O => \N__37264\,
            I => \N__37253\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__37259\,
            I => \N__37248\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37248\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__37253\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__37248\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37243\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37237\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__37234\,
            I => \N__37231\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37228\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37225\
        );

    \I__7622\ : Span4Mux_v
    port map (
            O => \N__37225\,
            I => \N__37220\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37217\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37214\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__37220\,
            I => \N__37211\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37208\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37204\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__37211\,
            I => \N__37201\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__37208\,
            I => \N__37198\
        );

    \I__7614\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37195\
        );

    \I__7613\ : Span4Mux_v
    port map (
            O => \N__37204\,
            I => \N__37190\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__37201\,
            I => \N__37190\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__37198\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37195\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__37190\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__7608\ : InMux
    port map (
            O => \N__37183\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37180\,
            I => \N__37177\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37177\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__37174\,
            I => \N__37171\
        );

    \I__7604\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37167\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__37170\,
            I => \N__37164\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__37167\,
            I => \N__37160\
        );

    \I__7601\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37157\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37154\
        );

    \I__7599\ : Sp12to4
    port map (
            O => \N__37160\,
            I => \N__37150\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37145\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37154\,
            I => \N__37145\
        );

    \I__7596\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37142\
        );

    \I__7595\ : Span12Mux_v
    port map (
            O => \N__37150\,
            I => \N__37139\
        );

    \I__7594\ : Span4Mux_v
    port map (
            O => \N__37145\,
            I => \N__37136\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__37142\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7592\ : Odrv12
    port map (
            O => \N__37139\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__37136\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37129\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37126\,
            I => \N__37121\
        );

    \I__7588\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37116\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37116\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37110\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37110\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__37115\,
            I => \N__37107\
        );

    \I__7583\ : Sp12to4
    port map (
            O => \N__37110\,
            I => \N__37104\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37101\
        );

    \I__7581\ : Span12Mux_v
    port map (
            O => \N__37104\,
            I => \N__37098\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37101\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7579\ : Odrv12
    port map (
            O => \N__37098\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37090\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__37090\,
            I => \N__37087\
        );

    \I__7576\ : Odrv12
    port map (
            O => \N__37087\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__37084\,
            I => \N__37081\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37077\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37080\,
            I => \N__37074\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__37077\,
            I => \N__37071\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37074\,
            I => \N__37068\
        );

    \I__7570\ : Sp12to4
    port map (
            O => \N__37071\,
            I => \N__37065\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__37068\,
            I => \N__37061\
        );

    \I__7568\ : Span12Mux_v
    port map (
            O => \N__37065\,
            I => \N__37058\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37055\
        );

    \I__7566\ : Sp12to4
    port map (
            O => \N__37061\,
            I => \N__37050\
        );

    \I__7565\ : Span12Mux_h
    port map (
            O => \N__37058\,
            I => \N__37050\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__37055\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__7563\ : Odrv12
    port map (
            O => \N__37050\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37045\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__7561\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37039\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37039\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__7559\ : CascadeMux
    port map (
            O => \N__37036\,
            I => \N__37032\
        );

    \I__7558\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37029\
        );

    \I__7557\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37026\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__37029\,
            I => \N__37022\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__37026\,
            I => \N__37019\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37016\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__37022\,
            I => \N__37013\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__37019\,
            I => \N__37010\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37007\
        );

    \I__7550\ : Sp12to4
    port map (
            O => \N__37013\,
            I => \N__37001\
        );

    \I__7549\ : Sp12to4
    port map (
            O => \N__37010\,
            I => \N__37001\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__37007\,
            I => \N__36998\
        );

    \I__7547\ : InMux
    port map (
            O => \N__37006\,
            I => \N__36995\
        );

    \I__7546\ : Span12Mux_h
    port map (
            O => \N__37001\,
            I => \N__36992\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__36998\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__36995\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__7543\ : Odrv12
    port map (
            O => \N__36992\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36985\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__7541\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__36979\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__36976\,
            I => \N__36972\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36975\,
            I => \N__36969\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36966\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36969\,
            I => \N__36962\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36966\,
            I => \N__36959\
        );

    \I__7534\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36956\
        );

    \I__7533\ : Span4Mux_v
    port map (
            O => \N__36962\,
            I => \N__36953\
        );

    \I__7532\ : Span4Mux_v
    port map (
            O => \N__36959\,
            I => \N__36950\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__36956\,
            I => \N__36947\
        );

    \I__7530\ : Sp12to4
    port map (
            O => \N__36953\,
            I => \N__36941\
        );

    \I__7529\ : Sp12to4
    port map (
            O => \N__36950\,
            I => \N__36941\
        );

    \I__7528\ : Span4Mux_v
    port map (
            O => \N__36947\,
            I => \N__36938\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36935\
        );

    \I__7526\ : Span12Mux_h
    port map (
            O => \N__36941\,
            I => \N__36932\
        );

    \I__7525\ : Odrv4
    port map (
            O => \N__36938\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36935\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__7523\ : Odrv12
    port map (
            O => \N__36932\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36925\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36922\,
            I => \N__36919\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36916\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36916\,
            I => \N__36911\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36907\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36904\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__36911\,
            I => \N__36901\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36898\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36907\,
            I => \N__36895\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__36904\,
            I => \N__36892\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__36901\,
            I => \N__36889\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36898\,
            I => \N__36886\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__36895\,
            I => \N__36883\
        );

    \I__7509\ : Span4Mux_h
    port map (
            O => \N__36892\,
            I => \N__36880\
        );

    \I__7508\ : Sp12to4
    port map (
            O => \N__36889\,
            I => \N__36877\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__36886\,
            I => \N__36874\
        );

    \I__7506\ : Odrv4
    port map (
            O => \N__36883\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__36880\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__7504\ : Odrv12
    port map (
            O => \N__36877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__36874\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36865\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36859\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36859\,
            I => \N__36856\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__36856\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__7498\ : CascadeMux
    port map (
            O => \N__36853\,
            I => \N__36850\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36845\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36842\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__36848\,
            I => \N__36839\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36836\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36833\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36839\,
            I => \N__36830\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__36836\,
            I => \N__36827\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__36833\,
            I => \N__36824\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__36830\,
            I => \N__36821\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__36827\,
            I => \N__36817\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__36824\,
            I => \N__36814\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__36821\,
            I => \N__36811\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36808\
        );

    \I__7484\ : Sp12to4
    port map (
            O => \N__36817\,
            I => \N__36805\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__36814\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__36811\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36808\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7480\ : Odrv12
    port map (
            O => \N__36805\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36796\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36793\,
            I => \N__36787\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36787\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36787\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__36784\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36775\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36775\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__36775\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36768\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36764\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36768\,
            I => \N__36761\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36767\,
            I => \N__36758\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36764\,
            I => \N__36755\
        );

    \I__7466\ : Span4Mux_v
    port map (
            O => \N__36761\,
            I => \N__36750\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36750\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__36755\,
            I => \N__36747\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__36750\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__36747\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36738\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36735\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__36738\,
            I => \N__36732\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36729\
        );

    \I__7457\ : Span4Mux_s3_h
    port map (
            O => \N__36732\,
            I => \N__36726\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__36729\,
            I => \N__36723\
        );

    \I__7455\ : Span4Mux_h
    port map (
            O => \N__36726\,
            I => \N__36720\
        );

    \I__7454\ : Odrv4
    port map (
            O => \N__36723\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__36720\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36711\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36708\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__36711\,
            I => \N__36705\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36708\,
            I => \N__36702\
        );

    \I__7448\ : Span4Mux_h
    port map (
            O => \N__36705\,
            I => \N__36699\
        );

    \I__7447\ : Span4Mux_s3_h
    port map (
            O => \N__36702\,
            I => \N__36696\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__36699\,
            I => \N__36693\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__36696\,
            I => \N__36690\
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__36693\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36690\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36685\,
            I => \N__36681\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36678\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36675\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36672\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__36675\,
            I => \N__36669\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__36672\,
            I => \N__36666\
        );

    \I__7436\ : Sp12to4
    port map (
            O => \N__36669\,
            I => \N__36663\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__36666\,
            I => \N__36660\
        );

    \I__7434\ : Odrv12
    port map (
            O => \N__36663\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__36660\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36649\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36649\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36649\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36642\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36639\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36642\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__36639\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36630\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36627\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36630\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__36627\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__7421\ : CascadeMux
    port map (
            O => \N__36622\,
            I => \N__36619\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36619\,
            I => \N__36616\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__36616\,
            I => \N__36613\
        );

    \I__7418\ : Odrv4
    port map (
            O => \N__36613\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__7417\ : CascadeMux
    port map (
            O => \N__36610\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36604\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36604\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\
        );

    \I__7414\ : CascadeMux
    port map (
            O => \N__36601\,
            I => \N__36597\
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__36600\,
            I => \N__36594\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36589\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36589\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36589\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__7409\ : CascadeMux
    port map (
            O => \N__36586\,
            I => \N__36583\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36583\,
            I => \N__36578\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36582\,
            I => \N__36575\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36572\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36578\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__36575\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__36572\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36565\,
            I => \bfn_14_10_0_\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__36562\,
            I => \N__36559\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36554\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36551\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36548\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__36554\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__36551\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36548\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36541\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36534\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36531\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__36534\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36531\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__36526\,
            I => \N__36523\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36518\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36515\
        );

    \I__7386\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36512\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__36518\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36515\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__36512\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36505\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36498\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36495\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36498\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36495\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__36490\,
            I => \N__36487\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36482\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36479\
        );

    \I__7374\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36476\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36482\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__36479\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__36476\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36469\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36466\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7368\ : CEMux
    port map (
            O => \N__36463\,
            I => \N__36457\
        );

    \I__7367\ : CEMux
    port map (
            O => \N__36462\,
            I => \N__36454\
        );

    \I__7366\ : CEMux
    port map (
            O => \N__36461\,
            I => \N__36451\
        );

    \I__7365\ : CEMux
    port map (
            O => \N__36460\,
            I => \N__36448\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N__36444\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__36454\,
            I => \N__36441\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36438\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36448\,
            I => \N__36435\
        );

    \I__7360\ : CEMux
    port map (
            O => \N__36447\,
            I => \N__36432\
        );

    \I__7359\ : Span4Mux_h
    port map (
            O => \N__36444\,
            I => \N__36429\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36426\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__36438\,
            I => \N__36423\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__36435\,
            I => \N__36420\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__36432\,
            I => \N__36417\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__36429\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__36426\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7352\ : Odrv4
    port map (
            O => \N__36423\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__36420\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7350\ : Odrv12
    port map (
            O => \N__36417\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7349\ : CascadeMux
    port map (
            O => \N__36406\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__36403\,
            I => \N__36400\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36394\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36394\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__36394\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__7344\ : CascadeMux
    port map (
            O => \N__36391\,
            I => \N__36388\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36383\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36380\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36386\,
            I => \N__36377\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36383\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__36380\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__36377\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36370\,
            I => \bfn_14_9_0_\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__36367\,
            I => \N__36364\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36359\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36356\
        );

    \I__7333\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36353\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36359\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__36356\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36353\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__7329\ : InMux
    port map (
            O => \N__36346\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36338\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36333\
        );

    \I__7326\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36333\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36338\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36333\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__7323\ : InMux
    port map (
            O => \N__36328\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__36325\,
            I => \N__36322\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36317\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36314\
        );

    \I__7319\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36311\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36314\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__36311\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36304\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__36301\,
            I => \N__36296\
        );

    \I__7313\ : CascadeMux
    port map (
            O => \N__36300\,
            I => \N__36293\
        );

    \I__7312\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36290\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36285\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36285\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36290\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__36285\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36280\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__36277\,
            I => \N__36274\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36269\
        );

    \I__7304\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36266\
        );

    \I__7303\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36263\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36269\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__36266\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36263\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36256\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7298\ : CascadeMux
    port map (
            O => \N__36253\,
            I => \N__36250\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36245\
        );

    \I__7296\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36242\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36239\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__36245\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36242\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36239\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36232\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__36229\,
            I => \N__36226\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36221\
        );

    \I__7288\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36218\
        );

    \I__7287\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36215\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__36221\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__36218\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36215\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36208\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7282\ : InMux
    port map (
            O => \N__36205\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__36202\,
            I => \N__36199\
        );

    \I__7280\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36194\
        );

    \I__7279\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36191\
        );

    \I__7278\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36188\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__36194\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__36191\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__36188\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__7274\ : InMux
    port map (
            O => \N__36181\,
            I => \bfn_14_8_0_\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__36178\,
            I => \N__36175\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36170\
        );

    \I__7271\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36167\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36164\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36170\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__36167\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36164\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36157\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__36154\,
            I => \N__36151\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36146\
        );

    \I__7263\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36143\
        );

    \I__7262\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36140\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__36146\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36143\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__36140\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36133\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__36130\,
            I => \N__36127\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36127\,
            I => \N__36122\
        );

    \I__7255\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36119\
        );

    \I__7254\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36116\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__36122\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__36119\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36116\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36109\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7249\ : CascadeMux
    port map (
            O => \N__36106\,
            I => \N__36103\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36098\
        );

    \I__7247\ : InMux
    port map (
            O => \N__36102\,
            I => \N__36095\
        );

    \I__7246\ : InMux
    port map (
            O => \N__36101\,
            I => \N__36092\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__36098\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__36095\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__36092\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36085\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__36082\,
            I => \N__36079\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36074\
        );

    \I__7239\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36071\
        );

    \I__7238\ : InMux
    port map (
            O => \N__36077\,
            I => \N__36068\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__36074\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__36071\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__36068\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36061\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__36058\,
            I => \N__36055\
        );

    \I__7232\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36050\
        );

    \I__7231\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36047\
        );

    \I__7230\ : InMux
    port map (
            O => \N__36053\,
            I => \N__36044\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__36050\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__36047\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__36044\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36037\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__36034\,
            I => \N__36031\
        );

    \I__7224\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36026\
        );

    \I__7223\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36023\
        );

    \I__7222\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36020\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__36026\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36023\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__36020\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__7218\ : InMux
    port map (
            O => \N__36013\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__36010\,
            I => \N__36006\
        );

    \I__7216\ : InMux
    port map (
            O => \N__36009\,
            I => \N__36002\
        );

    \I__7215\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35999\
        );

    \I__7214\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35996\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__36002\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35999\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__35996\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__35989\,
            I => \N__35985\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35981\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35978\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35975\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__35981\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35978\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__35975\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__7203\ : InMux
    port map (
            O => \N__35968\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__35965\,
            I => \N__35962\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35957\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35954\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35951\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35957\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__35954\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__35951\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35944\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35933\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35930\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35927\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35933\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35930\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__35927\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35920\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__35917\,
            I => \N__35914\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35909\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35906\
        );

    \I__7183\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35903\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__35909\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__35906\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35903\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__7179\ : InMux
    port map (
            O => \N__35896\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7178\ : CascadeMux
    port map (
            O => \N__35893\,
            I => \N__35890\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35885\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35882\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35879\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__35885\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__35882\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35879\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35872\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__35869\,
            I => \N__35866\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35861\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35858\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35855\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__35861\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35858\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__35855\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35848\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7162\ : CascadeMux
    port map (
            O => \N__35845\,
            I => \N__35842\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35842\,
            I => \N__35837\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35834\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35831\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__35837\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35834\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__35831\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35824\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35821\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35818\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35815\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35812\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__7150\ : InMux
    port map (
            O => \N__35809\,
            I => \bfn_13_27_0_\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35806\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__7148\ : CascadeMux
    port map (
            O => \N__35803\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\
        );

    \I__7147\ : CascadeMux
    port map (
            O => \N__35800\,
            I => \N__35797\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35794\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35794\,
            I => \N__35791\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35791\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35783\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35780\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35777\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35783\,
            I => \N__35774\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35780\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35777\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35774\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35764\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__35764\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35756\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35760\,
            I => \N__35753\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35750\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__35756\,
            I => \N__35747\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35753\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35750\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__35747\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35737\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35737\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35729\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35726\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35723\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35729\,
            I => \N__35718\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35726\,
            I => \N__35718\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35723\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__35718\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35710\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__7116\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35702\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35699\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35696\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35702\,
            I => \N__35693\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35699\,
            I => \N__35690\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35696\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__35693\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__35690\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35680\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__35680\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35677\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__7105\ : IoInMux
    port map (
            O => \N__35674\,
            I => \N__35671\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__35671\,
            I => \N__35668\
        );

    \I__7103\ : IoSpan4Mux
    port map (
            O => \N__35668\,
            I => \N__35665\
        );

    \I__7102\ : Sp12to4
    port map (
            O => \N__35665\,
            I => \N__35662\
        );

    \I__7101\ : Span12Mux_s10_v
    port map (
            O => \N__35662\,
            I => \N__35659\
        );

    \I__7100\ : Span12Mux_v
    port map (
            O => \N__35659\,
            I => \N__35656\
        );

    \I__7099\ : Span12Mux_h
    port map (
            O => \N__35656\,
            I => \N__35653\
        );

    \I__7098\ : Odrv12
    port map (
            O => \N__35653\,
            I => pwm_output_c
        );

    \I__7097\ : InMux
    port map (
            O => \N__35650\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35647\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35640\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35637\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35640\,
            I => \N__35634\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35637\,
            I => \N__35631\
        );

    \I__7091\ : Span4Mux_s3_h
    port map (
            O => \N__35634\,
            I => \N__35628\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__35631\,
            I => \N__35625\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__35628\,
            I => \N__35622\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__35625\,
            I => \N__35619\
        );

    \I__7087\ : Sp12to4
    port map (
            O => \N__35622\,
            I => \N__35616\
        );

    \I__7086\ : Odrv4
    port map (
            O => \N__35619\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__7085\ : Odrv12
    port map (
            O => \N__35616\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35596\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35596\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35584\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35584\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35584\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35584\
        );

    \I__7078\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35584\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35557\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35557\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35554\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35548\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35545\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35531\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35528\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35525\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35520\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35520\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35513\
        );

    \I__7066\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35513\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35513\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35502\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35502\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35502\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35502\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35502\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35572\,
            I => \N__35493\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35486\
        );

    \I__7057\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35486\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35486\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35471\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35471\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35471\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35471\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35471\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35471\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35471\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__35557\,
            I => \N__35468\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__35554\,
            I => \N__35465\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35460\
        );

    \I__7045\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35460\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35457\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35444\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__35545\,
            I => \N__35444\
        );

    \I__7041\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35431\
        );

    \I__7040\ : InMux
    port map (
            O => \N__35543\,
            I => \N__35431\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35431\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35431\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35431\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35431\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35415\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35415\
        );

    \I__7033\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35415\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35412\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35409\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35396\
        );

    \I__7029\ : Span4Mux_v
    port map (
            O => \N__35528\,
            I => \N__35396\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__35525\,
            I => \N__35396\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35396\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35513\,
            I => \N__35396\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35502\,
            I => \N__35396\
        );

    \I__7024\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35383\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35383\
        );

    \I__7022\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35383\
        );

    \I__7021\ : InMux
    port map (
            O => \N__35498\,
            I => \N__35383\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35383\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35383\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35493\,
            I => \N__35374\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35486\,
            I => \N__35374\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35374\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__35468\,
            I => \N__35374\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__35465\,
            I => \N__35369\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35369\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__35457\,
            I => \N__35366\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35349\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35455\,
            I => \N__35349\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35349\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35349\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35349\
        );

    \I__7006\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35349\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35349\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35349\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__35444\,
            I => \N__35344\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35344\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35331\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35331\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35331\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35331\
        );

    \I__6997\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35331\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35331\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35324\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35324\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35324\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35415\,
            I => \N__35321\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35412\,
            I => \N__35314\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35409\,
            I => \N__35314\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__35396\,
            I => \N__35314\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35307\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__35374\,
            I => \N__35307\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__35369\,
            I => \N__35307\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__35366\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__35349\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__35344\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35331\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35324\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6980\ : Odrv12
    port map (
            O => \N__35321\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6979\ : Odrv4
    port map (
            O => \N__35314\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6978\ : Odrv4
    port map (
            O => \N__35307\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6977\ : CascadeMux
    port map (
            O => \N__35290\,
            I => \N__35287\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35284\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__35284\,
            I => \N__35280\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35276\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__35280\,
            I => \N__35273\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35270\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35267\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__35273\,
            I => \N__35263\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35260\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__35267\,
            I => \N__35257\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35266\,
            I => \N__35254\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__35263\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6965\ : Odrv12
    port map (
            O => \N__35260\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6964\ : Odrv4
    port map (
            O => \N__35257\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__35254\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35210\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35244\,
            I => \N__35210\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35199\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35199\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35199\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35199\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35199\
        );

    \I__6955\ : CascadeMux
    port map (
            O => \N__35238\,
            I => \N__35194\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35189\
        );

    \I__6953\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35181\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__35235\,
            I => \N__35178\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__35234\,
            I => \N__35172\
        );

    \I__6950\ : CascadeMux
    port map (
            O => \N__35233\,
            I => \N__35168\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__35232\,
            I => \N__35165\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35150\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35150\
        );

    \I__6946\ : InMux
    port map (
            O => \N__35229\,
            I => \N__35150\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35150\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35150\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35150\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__35225\,
            I => \N__35128\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__35224\,
            I => \N__35124\
        );

    \I__6940\ : CascadeMux
    port map (
            O => \N__35223\,
            I => \N__35120\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__35222\,
            I => \N__35116\
        );

    \I__6938\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35093\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35093\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35093\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35093\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35093\
        );

    \I__6933\ : InMux
    port map (
            O => \N__35216\,
            I => \N__35093\
        );

    \I__6932\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35093\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__35210\,
            I => \N__35088\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__35199\,
            I => \N__35088\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35198\,
            I => \N__35085\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35080\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35080\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__35193\,
            I => \N__35077\
        );

    \I__6925\ : CascadeMux
    port map (
            O => \N__35192\,
            I => \N__35073\
        );

    \I__6924\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35069\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35062\
        );

    \I__6922\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35062\
        );

    \I__6921\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35062\
        );

    \I__6920\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35057\
        );

    \I__6919\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35057\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35181\,
            I => \N__35054\
        );

    \I__6917\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35051\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35038\
        );

    \I__6915\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35038\
        );

    \I__6914\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35038\
        );

    \I__6913\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35038\
        );

    \I__6912\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35038\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35038\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35031\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35031\
        );

    \I__6908\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35031\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35150\,
            I => \N__35028\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35023\
        );

    \I__6905\ : InMux
    port map (
            O => \N__35148\,
            I => \N__35023\
        );

    \I__6904\ : CascadeMux
    port map (
            O => \N__35147\,
            I => \N__35020\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__35146\,
            I => \N__35017\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__35145\,
            I => \N__35009\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__35144\,
            I => \N__35005\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__35143\,
            I => \N__35001\
        );

    \I__6899\ : InMux
    port map (
            O => \N__35142\,
            I => \N__34993\
        );

    \I__6898\ : InMux
    port map (
            O => \N__35141\,
            I => \N__34993\
        );

    \I__6897\ : InMux
    port map (
            O => \N__35140\,
            I => \N__34993\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__35139\,
            I => \N__34990\
        );

    \I__6895\ : CascadeMux
    port map (
            O => \N__35138\,
            I => \N__34986\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__35137\,
            I => \N__34982\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__35136\,
            I => \N__34978\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35135\,
            I => \N__34966\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35134\,
            I => \N__34966\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35133\,
            I => \N__34966\
        );

    \I__6889\ : InMux
    port map (
            O => \N__35132\,
            I => \N__34966\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35131\,
            I => \N__34966\
        );

    \I__6887\ : InMux
    port map (
            O => \N__35128\,
            I => \N__34949\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35127\,
            I => \N__34949\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35124\,
            I => \N__34949\
        );

    \I__6884\ : InMux
    port map (
            O => \N__35123\,
            I => \N__34949\
        );

    \I__6883\ : InMux
    port map (
            O => \N__35120\,
            I => \N__34949\
        );

    \I__6882\ : InMux
    port map (
            O => \N__35119\,
            I => \N__34949\
        );

    \I__6881\ : InMux
    port map (
            O => \N__35116\,
            I => \N__34949\
        );

    \I__6880\ : InMux
    port map (
            O => \N__35115\,
            I => \N__34949\
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__35114\,
            I => \N__34946\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__35113\,
            I => \N__34942\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__35112\,
            I => \N__34938\
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__35111\,
            I => \N__34934\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__35110\,
            I => \N__34930\
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__35109\,
            I => \N__34926\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__35108\,
            I => \N__34922\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__34918\
        );

    \I__6871\ : Span4Mux_h
    port map (
            O => \N__35088\,
            I => \N__34911\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__35085\,
            I => \N__34911\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__35080\,
            I => \N__34911\
        );

    \I__6868\ : InMux
    port map (
            O => \N__35077\,
            I => \N__34908\
        );

    \I__6867\ : InMux
    port map (
            O => \N__35076\,
            I => \N__34903\
        );

    \I__6866\ : InMux
    port map (
            O => \N__35073\,
            I => \N__34903\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__35072\,
            I => \N__34897\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35069\,
            I => \N__34890\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__34885\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35057\,
            I => \N__34885\
        );

    \I__6861\ : Span4Mux_v
    port map (
            O => \N__35054\,
            I => \N__34876\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__35051\,
            I => \N__34876\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__34876\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__34876\
        );

    \I__6857\ : Span4Mux_h
    port map (
            O => \N__35028\,
            I => \N__34864\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__34864\
        );

    \I__6855\ : InMux
    port map (
            O => \N__35020\,
            I => \N__34851\
        );

    \I__6854\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34851\
        );

    \I__6853\ : InMux
    port map (
            O => \N__35016\,
            I => \N__34851\
        );

    \I__6852\ : InMux
    port map (
            O => \N__35015\,
            I => \N__34851\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35014\,
            I => \N__34851\
        );

    \I__6850\ : InMux
    port map (
            O => \N__35013\,
            I => \N__34851\
        );

    \I__6849\ : InMux
    port map (
            O => \N__35012\,
            I => \N__34836\
        );

    \I__6848\ : InMux
    port map (
            O => \N__35009\,
            I => \N__34836\
        );

    \I__6847\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34836\
        );

    \I__6846\ : InMux
    port map (
            O => \N__35005\,
            I => \N__34836\
        );

    \I__6845\ : InMux
    port map (
            O => \N__35004\,
            I => \N__34836\
        );

    \I__6844\ : InMux
    port map (
            O => \N__35001\,
            I => \N__34836\
        );

    \I__6843\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34836\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34993\,
            I => \N__34833\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34816\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34816\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34816\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34816\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34816\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34816\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34816\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34816\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34811\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34811\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34794\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34794\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34794\
        );

    \I__6828\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34794\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34794\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34794\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34794\
        );

    \I__6824\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34794\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34781\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34781\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34781\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34781\
        );

    \I__6819\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34781\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34781\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__34918\,
            I => \N__34772\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__34911\,
            I => \N__34772\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34772\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__34903\,
            I => \N__34772\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34755\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34755\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34755\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34755\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34755\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34755\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34755\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34755\
        );

    \I__6805\ : Span4Mux_h
    port map (
            O => \N__34890\,
            I => \N__34750\
        );

    \I__6804\ : Span4Mux_h
    port map (
            O => \N__34885\,
            I => \N__34750\
        );

    \I__6803\ : Span4Mux_v
    port map (
            O => \N__34876\,
            I => \N__34747\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__34875\,
            I => \N__34744\
        );

    \I__6801\ : CascadeMux
    port map (
            O => \N__34874\,
            I => \N__34740\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__34873\,
            I => \N__34736\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__34872\,
            I => \N__34732\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__34871\,
            I => \N__34728\
        );

    \I__6797\ : CascadeMux
    port map (
            O => \N__34870\,
            I => \N__34724\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__34869\,
            I => \N__34720\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__34864\,
            I => \N__34702\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34702\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N__34702\
        );

    \I__6792\ : Span4Mux_v
    port map (
            O => \N__34833\,
            I => \N__34702\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34702\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__34811\,
            I => \N__34702\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34702\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__34781\,
            I => \N__34702\
        );

    \I__6787\ : Span4Mux_v
    port map (
            O => \N__34772\,
            I => \N__34699\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34696\
        );

    \I__6785\ : Span4Mux_v
    port map (
            O => \N__34750\,
            I => \N__34691\
        );

    \I__6784\ : Span4Mux_v
    port map (
            O => \N__34747\,
            I => \N__34691\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34674\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34674\
        );

    \I__6781\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34674\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34674\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34674\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34674\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34732\,
            I => \N__34674\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34731\,
            I => \N__34674\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34661\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34661\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34661\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34661\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34720\,
            I => \N__34661\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34661\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__34702\,
            I => \N__34658\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__34699\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__34696\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6766\ : Odrv4
    port map (
            O => \N__34691\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34674\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34661\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6763\ : Odrv4
    port map (
            O => \N__34658\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34642\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34642\,
            I => \N__34639\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__34639\,
            I => \N__34634\
        );

    \I__6759\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34631\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34628\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__34634\,
            I => \N__34623\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34631\,
            I => \N__34623\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34620\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__34623\,
            I => \N__34617\
        );

    \I__6753\ : Span12Mux_s11_h
    port map (
            O => \N__34620\,
            I => \N__34614\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__34617\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__6751\ : Odrv12
    port map (
            O => \N__34614\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34606\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34603\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__34603\,
            I => \N__34600\
        );

    \I__6747\ : Odrv4
    port map (
            O => \N__34600\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34594\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34589\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34586\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34583\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__34589\,
            I => \N__34580\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34577\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34583\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6739\ : Odrv4
    port map (
            O => \N__34580\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__34577\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__34567\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34560\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34557\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__34560\,
            I => \N__34551\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__34557\,
            I => \N__34551\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34548\
        );

    \I__6730\ : Span4Mux_h
    port map (
            O => \N__34551\,
            I => \N__34545\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34548\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__6728\ : Odrv4
    port map (
            O => \N__34545\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__34540\,
            I => \N__34537\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34534\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__34534\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34528\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__34528\,
            I => \N__34523\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34520\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34517\
        );

    \I__6720\ : Span4Mux_v
    port map (
            O => \N__34523\,
            I => \N__34514\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__34520\,
            I => \N__34511\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__34517\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__34514\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__34511\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__34504\,
            I => \N__34501\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34498\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34498\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34490\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34487\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34484\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34490\,
            I => \N__34479\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34487\,
            I => \N__34479\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__34484\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__34479\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__6705\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34471\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__34471\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34463\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34460\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34457\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34463\,
            I => \N__34452\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34460\,
            I => \N__34452\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__34457\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__34452\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__34447\,
            I => \N__34444\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34441\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34438\,
            I => \N__34433\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34430\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34427\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34424\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__34430\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__34427\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__34424\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34414\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34414\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34408\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__34408\,
            I => \N__34404\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34401\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__34404\,
            I => \N__34398\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34395\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__34398\,
            I => \N__34392\
        );

    \I__6678\ : Span12Mux_s7_h
    port map (
            O => \N__34395\,
            I => \N__34389\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__34392\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6676\ : Odrv12
    port map (
            O => \N__34389\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34380\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34377\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34374\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34371\
        );

    \I__6671\ : Span4Mux_h
    port map (
            O => \N__34374\,
            I => \N__34368\
        );

    \I__6670\ : Span4Mux_s3_h
    port map (
            O => \N__34371\,
            I => \N__34365\
        );

    \I__6669\ : Span4Mux_h
    port map (
            O => \N__34368\,
            I => \N__34362\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__34365\,
            I => \N__34359\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__34362\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__34359\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34350\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34353\,
            I => \N__34347\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__34350\,
            I => \N__34344\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__34347\,
            I => \N__34341\
        );

    \I__6661\ : Sp12to4
    port map (
            O => \N__34344\,
            I => \N__34338\
        );

    \I__6660\ : Span12Mux_v
    port map (
            O => \N__34341\,
            I => \N__34333\
        );

    \I__6659\ : Span12Mux_v
    port map (
            O => \N__34338\,
            I => \N__34333\
        );

    \I__6658\ : Odrv12
    port map (
            O => \N__34333\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34326\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34323\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34326\,
            I => \N__34320\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__34323\,
            I => \N__34317\
        );

    \I__6653\ : Span4Mux_s3_h
    port map (
            O => \N__34320\,
            I => \N__34314\
        );

    \I__6652\ : Span4Mux_v
    port map (
            O => \N__34317\,
            I => \N__34311\
        );

    \I__6651\ : Sp12to4
    port map (
            O => \N__34314\,
            I => \N__34308\
        );

    \I__6650\ : Sp12to4
    port map (
            O => \N__34311\,
            I => \N__34303\
        );

    \I__6649\ : Span12Mux_v
    port map (
            O => \N__34308\,
            I => \N__34303\
        );

    \I__6648\ : Odrv12
    port map (
            O => \N__34303\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34296\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34293\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34290\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__34293\,
            I => \N__34287\
        );

    \I__6643\ : Span4Mux_v
    port map (
            O => \N__34290\,
            I => \N__34284\
        );

    \I__6642\ : Span4Mux_v
    port map (
            O => \N__34287\,
            I => \N__34281\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__34284\,
            I => \N__34276\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__34281\,
            I => \N__34276\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__34276\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34269\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34272\,
            I => \N__34266\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34263\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34260\
        );

    \I__6634\ : Span4Mux_s2_h
    port map (
            O => \N__34263\,
            I => \N__34257\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__34260\,
            I => \N__34254\
        );

    \I__6632\ : Sp12to4
    port map (
            O => \N__34257\,
            I => \N__34251\
        );

    \I__6631\ : Sp12to4
    port map (
            O => \N__34254\,
            I => \N__34246\
        );

    \I__6630\ : Span12Mux_v
    port map (
            O => \N__34251\,
            I => \N__34246\
        );

    \I__6629\ : Odrv12
    port map (
            O => \N__34246\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34239\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34236\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__34239\,
            I => \N__34233\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34236\,
            I => \N__34230\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__34233\,
            I => \N__34227\
        );

    \I__6623\ : Span4Mux_h
    port map (
            O => \N__34230\,
            I => \N__34224\
        );

    \I__6622\ : Sp12to4
    port map (
            O => \N__34227\,
            I => \N__34221\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__34224\,
            I => \N__34218\
        );

    \I__6620\ : Span12Mux_s7_h
    port map (
            O => \N__34221\,
            I => \N__34215\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__34218\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__6618\ : Odrv12
    port map (
            O => \N__34215\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__6617\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34206\
        );

    \I__6616\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34203\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__34206\,
            I => \N__34200\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34197\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__34200\,
            I => \N__34194\
        );

    \I__6612\ : Span4Mux_h
    port map (
            O => \N__34197\,
            I => \N__34191\
        );

    \I__6611\ : Sp12to4
    port map (
            O => \N__34194\,
            I => \N__34188\
        );

    \I__6610\ : Span4Mux_h
    port map (
            O => \N__34191\,
            I => \N__34185\
        );

    \I__6609\ : Span12Mux_s7_h
    port map (
            O => \N__34188\,
            I => \N__34182\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__34185\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__6607\ : Odrv12
    port map (
            O => \N__34182\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34173\
        );

    \I__6605\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34170\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__34173\,
            I => \N__34167\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__34170\,
            I => \N__34164\
        );

    \I__6602\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__34161\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__34164\,
            I => \N__34158\
        );

    \I__6600\ : Sp12to4
    port map (
            O => \N__34161\,
            I => \N__34155\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__34158\,
            I => \N__34152\
        );

    \I__6598\ : Span12Mux_s7_h
    port map (
            O => \N__34155\,
            I => \N__34149\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__34152\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__6596\ : Odrv12
    port map (
            O => \N__34149\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__6595\ : IoInMux
    port map (
            O => \N__34144\,
            I => \N__34141\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34138\
        );

    \I__6593\ : Span12Mux_s10_v
    port map (
            O => \N__34138\,
            I => \N__34135\
        );

    \I__6592\ : Odrv12
    port map (
            O => \N__34135\,
            I => s2_phy_c
        );

    \I__6591\ : InMux
    port map (
            O => \N__34132\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34124\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34121\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34118\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34124\,
            I => \N__34115\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__34121\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__34118\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__34115\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34108\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34105\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__6580\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34094\
        );

    \I__6579\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34091\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34088\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34094\,
            I => \N__34085\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__34091\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34088\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6574\ : Odrv12
    port map (
            O => \N__34085\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__6573\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34074\
        );

    \I__6572\ : InMux
    port map (
            O => \N__34077\,
            I => \N__34071\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34074\,
            I => \N__34068\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34071\,
            I => \N__34065\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__34068\,
            I => \N__34062\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__34065\,
            I => \N__34059\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__34062\,
            I => \N__34056\
        );

    \I__6566\ : Sp12to4
    port map (
            O => \N__34059\,
            I => \N__34053\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__34056\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__6564\ : Odrv12
    port map (
            O => \N__34053\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34044\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34041\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34038\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__34035\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__34038\,
            I => \N__34032\
        );

    \I__6558\ : Span4Mux_s3_h
    port map (
            O => \N__34035\,
            I => \N__34029\
        );

    \I__6557\ : Span4Mux_h
    port map (
            O => \N__34032\,
            I => \N__34024\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__34029\,
            I => \N__34024\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__34024\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6554\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34018\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__34018\,
            I => \N__34015\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__34015\,
            I => \N__34011\
        );

    \I__6551\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34008\
        );

    \I__6550\ : Sp12to4
    port map (
            O => \N__34011\,
            I => \N__34005\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__34002\
        );

    \I__6548\ : Span12Mux_s7_h
    port map (
            O => \N__34005\,
            I => \N__33999\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__34002\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__6546\ : Odrv12
    port map (
            O => \N__33999\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33990\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33987\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33990\,
            I => \N__33984\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__33987\,
            I => \N__33981\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__33984\,
            I => \N__33978\
        );

    \I__6540\ : Span4Mux_v
    port map (
            O => \N__33981\,
            I => \N__33975\
        );

    \I__6539\ : Span4Mux_h
    port map (
            O => \N__33978\,
            I => \N__33972\
        );

    \I__6538\ : Span4Mux_h
    port map (
            O => \N__33975\,
            I => \N__33969\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__33972\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__33969\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33961\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33957\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33954\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__33957\,
            I => \N__33951\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__33954\,
            I => \N__33948\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__33951\,
            I => \N__33945\
        );

    \I__6529\ : Span12Mux_s7_h
    port map (
            O => \N__33948\,
            I => \N__33942\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__33945\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__6527\ : Odrv12
    port map (
            O => \N__33942\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33933\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33930\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33933\,
            I => \N__33927\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33924\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__33927\,
            I => \N__33921\
        );

    \I__6521\ : Span4Mux_v
    port map (
            O => \N__33924\,
            I => \N__33918\
        );

    \I__6520\ : Sp12to4
    port map (
            O => \N__33921\,
            I => \N__33915\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__33918\,
            I => \N__33912\
        );

    \I__6518\ : Span12Mux_s7_h
    port map (
            O => \N__33915\,
            I => \N__33909\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__33912\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__6516\ : Odrv12
    port map (
            O => \N__33909\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__6515\ : CascadeMux
    port map (
            O => \N__33904\,
            I => \N__33900\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33895\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33895\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33891\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33888\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__33891\,
            I => \N__33885\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__33888\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__33885\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33880\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__33877\,
            I => \N__33874\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33867\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33867\
        );

    \I__6503\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33864\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33867\,
            I => \N__33861\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__33864\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__33861\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33856\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33846\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33846\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33843\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33840\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33843\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__33840\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33835\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__33832\,
            I => \N__33829\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33823\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33823\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33823\,
            I => \N__33819\
        );

    \I__6487\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33816\
        );

    \I__6486\ : Span4Mux_h
    port map (
            O => \N__33819\,
            I => \N__33813\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33816\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__33813\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33808\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33798\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33798\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33795\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33792\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33795\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__33792\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33787\,
            I => \bfn_13_15_0_\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33779\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33774\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33774\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33779\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33774\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__6470\ : InMux
    port map (
            O => \N__33769\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__6469\ : CascadeMux
    port map (
            O => \N__33766\,
            I => \N__33762\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33758\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33762\,
            I => \N__33753\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33753\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__33758\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__33753\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33748\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__33745\,
            I => \N__33740\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33737\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33732\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33732\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__33737\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__33732\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33727\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33719\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33714\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33714\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33719\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__33714\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33705\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33702\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__33705\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33702\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33697\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33690\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33687\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33690\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33687\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33682\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33675\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33672\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33675\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33672\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33667\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33658\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33658\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__33658\,
            I => \N__33654\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33651\
        );

    \I__6431\ : Span4Mux_h
    port map (
            O => \N__33654\,
            I => \N__33648\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33651\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__33648\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33643\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__33640\,
            I => \N__33637\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33631\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33631\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33627\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33624\
        );

    \I__6422\ : Span4Mux_h
    port map (
            O => \N__33627\,
            I => \N__33621\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__33624\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__33621\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33616\,
            I => \bfn_13_14_0_\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__33613\,
            I => \N__33610\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33604\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33604\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33604\,
            I => \N__33600\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__33600\,
            I => \N__33594\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33597\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__33594\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33589\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33580\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33580\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33576\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33579\,
            I => \N__33573\
        );

    \I__6405\ : Span4Mux_h
    port map (
            O => \N__33576\,
            I => \N__33570\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__33573\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__33570\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33565\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33555\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33555\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33552\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33555\,
            I => \N__33549\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__33552\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__6396\ : Odrv4
    port map (
            O => \N__33549\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33544\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33537\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33540\,
            I => \N__33534\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33537\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__33534\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33529\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33522\
        );

    \I__6388\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33519\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__33522\,
            I => \N__33516\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__33519\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__33516\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33511\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33504\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33501\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__33504\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__33501\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33496\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33489\
        );

    \I__6377\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33486\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__33489\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33486\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6374\ : InMux
    port map (
            O => \N__33481\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33474\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33471\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33474\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__33471\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33466\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33459\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33456\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__33459\,
            I => \N__33453\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33456\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__33453\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6363\ : InMux
    port map (
            O => \N__33448\,
            I => \bfn_13_13_0_\
        );

    \I__6362\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33441\
        );

    \I__6361\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33438\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__33441\,
            I => \N__33435\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__33438\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__33435\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6357\ : InMux
    port map (
            O => \N__33430\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33423\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33426\,
            I => \N__33420\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__33423\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__33420\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33415\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33408\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33405\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__33408\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__33405\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33400\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33391\
        );

    \I__6345\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33391\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__33391\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33382\
        );

    \I__6342\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33382\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__33382\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33375\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33372\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33375\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__33372\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6336\ : InMux
    port map (
            O => \N__33367\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__33364\,
            I => \N__33361\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33357\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33354\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33357\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33354\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6330\ : InMux
    port map (
            O => \N__33349\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__6329\ : InMux
    port map (
            O => \N__33346\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33343\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33340\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33337\,
            I => \bfn_13_10_0_\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33334\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33331\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33328\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33325\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33284\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33284\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33284\
        );

    \I__6318\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33284\
        );

    \I__6317\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33275\
        );

    \I__6316\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33275\
        );

    \I__6315\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33275\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33275\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33268\
        );

    \I__6312\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33268\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33268\
        );

    \I__6310\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33259\
        );

    \I__6309\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33259\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33259\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33259\
        );

    \I__6306\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33252\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33252\
        );

    \I__6304\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33252\
        );

    \I__6303\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33243\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33243\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33243\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33243\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33234\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33234\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33234\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33234\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33225\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33225\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33225\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33225\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33220\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__33275\,
            I => \N__33220\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33215\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33259\,
            I => \N__33215\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33208\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33208\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__33234\,
            I => \N__33208\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33205\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__33220\,
            I => \N__33198\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__33215\,
            I => \N__33198\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__33208\,
            I => \N__33198\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__33205\,
            I => \N__33195\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__33198\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__33195\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6277\ : InMux
    port map (
            O => \N__33190\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6276\ : CEMux
    port map (
            O => \N__33187\,
            I => \N__33183\
        );

    \I__6275\ : CEMux
    port map (
            O => \N__33186\,
            I => \N__33178\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33175\
        );

    \I__6273\ : CEMux
    port map (
            O => \N__33182\,
            I => \N__33172\
        );

    \I__6272\ : CEMux
    port map (
            O => \N__33181\,
            I => \N__33169\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33178\,
            I => \N__33166\
        );

    \I__6270\ : Span4Mux_h
    port map (
            O => \N__33175\,
            I => \N__33163\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__33172\,
            I => \N__33160\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33169\,
            I => \N__33157\
        );

    \I__6267\ : Span4Mux_v
    port map (
            O => \N__33166\,
            I => \N__33154\
        );

    \I__6266\ : Span4Mux_v
    port map (
            O => \N__33163\,
            I => \N__33151\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33148\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__33157\,
            I => \N__33143\
        );

    \I__6263\ : Span4Mux_h
    port map (
            O => \N__33154\,
            I => \N__33143\
        );

    \I__6262\ : Odrv4
    port map (
            O => \N__33151\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__6261\ : Odrv4
    port map (
            O => \N__33148\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__33143\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33136\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6258\ : InMux
    port map (
            O => \N__33133\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33130\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33127\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33124\,
            I => \bfn_13_9_0_\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33121\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33118\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33115\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33112\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33109\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33106\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33103\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33100\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33097\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6245\ : InMux
    port map (
            O => \N__33094\,
            I => \bfn_13_8_0_\
        );

    \I__6244\ : InMux
    port map (
            O => \N__33091\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33088\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6242\ : InMux
    port map (
            O => \N__33085\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6241\ : InMux
    port map (
            O => \N__33082\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33079\,
            I => \bfn_12_27_0_\
        );

    \I__6239\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33062\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33062\
        );

    \I__6237\ : InMux
    port map (
            O => \N__33074\,
            I => \N__33053\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33073\,
            I => \N__33053\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33072\,
            I => \N__33053\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33071\,
            I => \N__33053\
        );

    \I__6233\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33044\
        );

    \I__6232\ : InMux
    port map (
            O => \N__33069\,
            I => \N__33044\
        );

    \I__6231\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33044\
        );

    \I__6230\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33044\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33041\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__33053\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__33044\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__33041\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33034\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__6224\ : IoInMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33025\
        );

    \I__6222\ : IoSpan4Mux
    port map (
            O => \N__33025\,
            I => \N__33022\
        );

    \I__6221\ : Span4Mux_s0_v
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__33019\,
            I => \GB_BUFFER_red_c_g_THRU_CO\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33016\,
            I => \bfn_13_7_0_\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33013\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__6217\ : InMux
    port map (
            O => \N__33010\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6216\ : InMux
    port map (
            O => \N__33007\,
            I => \N__33004\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__33004\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__33001\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32998\,
            I => \bfn_12_26_0_\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32995\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32992\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32989\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32986\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__6208\ : InMux
    port map (
            O => \N__32983\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32980\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__32971\,
            I => \N__32966\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32970\,
            I => \N__32963\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32960\
        );

    \I__6201\ : Odrv4
    port map (
            O => \N__32966\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__32963\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__32960\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32949\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32946\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32949\,
            I => \N__32941\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__32946\,
            I => \N__32941\
        );

    \I__6194\ : Span4Mux_h
    port map (
            O => \N__32941\,
            I => \N__32936\
        );

    \I__6193\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32931\
        );

    \I__6192\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32931\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__32936\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__32931\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__32926\,
            I => \N__32923\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__32917\,
            I => \N__32914\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__32914\,
            I => \N__32911\
        );

    \I__6184\ : Span4Mux_v
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__6183\ : Odrv4
    port map (
            O => \N__32908\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32902\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32902\,
            I => \N__32899\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__32899\,
            I => \N__32894\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32891\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32888\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__32894\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__32891\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32888\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6174\ : CEMux
    port map (
            O => \N__32881\,
            I => \N__32857\
        );

    \I__6173\ : CEMux
    port map (
            O => \N__32880\,
            I => \N__32857\
        );

    \I__6172\ : CEMux
    port map (
            O => \N__32879\,
            I => \N__32857\
        );

    \I__6171\ : CEMux
    port map (
            O => \N__32878\,
            I => \N__32857\
        );

    \I__6170\ : CEMux
    port map (
            O => \N__32877\,
            I => \N__32857\
        );

    \I__6169\ : CEMux
    port map (
            O => \N__32876\,
            I => \N__32857\
        );

    \I__6168\ : CEMux
    port map (
            O => \N__32875\,
            I => \N__32857\
        );

    \I__6167\ : CEMux
    port map (
            O => \N__32874\,
            I => \N__32857\
        );

    \I__6166\ : GlobalMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__6165\ : gio2CtrlBuf
    port map (
            O => \N__32854\,
            I => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32848\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32845\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__32845\,
            I => \N__32842\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__32842\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__6160\ : CascadeMux
    port map (
            O => \N__32839\,
            I => \N__32835\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32829\
        );

    \I__6158\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32829\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32826\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32823\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32826\,
            I => \N__32819\
        );

    \I__6154\ : Span12Mux_h
    port map (
            O => \N__32823\,
            I => \N__32816\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32813\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__32819\,
            I => \N__32810\
        );

    \I__6151\ : Odrv12
    port map (
            O => \N__32816\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__32813\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__32810\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__32803\,
            I => \N__32800\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32797\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32794\
        );

    \I__6145\ : Span4Mux_v
    port map (
            O => \N__32794\,
            I => \N__32791\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__32791\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32772\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32787\,
            I => \N__32769\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32764\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32764\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32748\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32748\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32748\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32748\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32748\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32748\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32745\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32740\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32735\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32775\,
            I => \N__32735\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32728\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32728\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32764\,
            I => \N__32728\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32721\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32721\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32721\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__32748\,
            I => \N__32718\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32745\,
            I => \N__32715\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32710\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32710\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32740\,
            I => \N__32705\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32735\,
            I => \N__32701\
        );

    \I__6117\ : Span4Mux_v
    port map (
            O => \N__32728\,
            I => \N__32690\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__32721\,
            I => \N__32690\
        );

    \I__6115\ : Span4Mux_h
    port map (
            O => \N__32718\,
            I => \N__32690\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__32715\,
            I => \N__32690\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32710\,
            I => \N__32690\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32685\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32685\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__32705\,
            I => \N__32679\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32676\
        );

    \I__6108\ : Span4Mux_v
    port map (
            O => \N__32701\,
            I => \N__32673\
        );

    \I__6107\ : Span4Mux_v
    port map (
            O => \N__32690\,
            I => \N__32668\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32685\,
            I => \N__32668\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32665\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32660\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32660\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__32679\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32676\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__32673\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6099\ : Odrv4
    port map (
            O => \N__32668\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__32665\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32660\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__32647\,
            I => \N__32644\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32635\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32635\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32635\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32635\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32620\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32620\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32620\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32620\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32620\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__32617\,
            I => \N__32614\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32611\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32608\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__32608\,
            I => \N__32605\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__32605\,
            I => \N__32602\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__32602\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__6080\ : CascadeMux
    port map (
            O => \N__32599\,
            I => \N__32593\
        );

    \I__6079\ : CascadeMux
    port map (
            O => \N__32598\,
            I => \N__32590\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32585\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32585\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32581\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32578\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32585\,
            I => \N__32575\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32572\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32581\,
            I => \N__32569\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__32578\,
            I => \N__32566\
        );

    \I__6070\ : Span4Mux_h
    port map (
            O => \N__32575\,
            I => \N__32563\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32560\
        );

    \I__6068\ : Span12Mux_s10_v
    port map (
            O => \N__32569\,
            I => \N__32557\
        );

    \I__6067\ : Span4Mux_h
    port map (
            O => \N__32566\,
            I => \N__32552\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__32563\,
            I => \N__32552\
        );

    \I__6065\ : Span4Mux_h
    port map (
            O => \N__32560\,
            I => \N__32549\
        );

    \I__6064\ : Odrv12
    port map (
            O => \N__32557\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__32552\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__32549\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32538\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32535\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32538\,
            I => \N__32529\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32535\,
            I => \N__32529\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32526\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__32529\,
            I => \N__32523\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32526\,
            I => \N__32520\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__32523\,
            I => \N__32517\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__32520\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__32517\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__32512\,
            I => \N__32509\
        );

    \I__6050\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32506\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32503\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__32503\,
            I => \N__32500\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__32500\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__32497\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__6045\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32491\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32485\
        );

    \I__6043\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32482\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32477\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32477\
        );

    \I__6040\ : Odrv12
    port map (
            O => \N__32485\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32482\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__32477\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__6037\ : CascadeMux
    port map (
            O => \N__32470\,
            I => \N__32466\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32463\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32459\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__32463\,
            I => \N__32456\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32453\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32459\,
            I => \N__32450\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__32456\,
            I => \N__32447\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__32453\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__32450\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__32447\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__6027\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32437\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32434\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__32434\,
            I => \N__32431\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__32431\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__32428\,
            I => \N__32425\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32421\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32418\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32415\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32412\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__32415\,
            I => \N__32408\
        );

    \I__6017\ : Sp12to4
    port map (
            O => \N__32412\,
            I => \N__32405\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32402\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__32408\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6014\ : Odrv12
    port map (
            O => \N__32405\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__32402\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__6012\ : CascadeMux
    port map (
            O => \N__32395\,
            I => \N__32392\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32388\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32385\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__32388\,
            I => \N__32382\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32377\
        );

    \I__6007\ : Span4Mux_v
    port map (
            O => \N__32382\,
            I => \N__32377\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__32377\,
            I => \N__32373\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32370\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__32373\,
            I => \N__32366\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32363\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32360\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__32366\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__32363\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__32360\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32350\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32350\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32344\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__32344\,
            I => \N__32341\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__32338\,
            I => \N__32335\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__32335\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32329\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__32329\,
            I => \N__32326\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__32326\,
            I => \N__32323\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__32323\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__5987\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32317\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32314\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__32314\,
            I => \N__32311\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__32311\,
            I => \N__32308\
        );

    \I__5983\ : Odrv4
    port map (
            O => \N__32308\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__5982\ : CascadeMux
    port map (
            O => \N__32305\,
            I => \N__32301\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32295\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32295\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32292\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32295\,
            I => \N__32287\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__32292\,
            I => \N__32287\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__32287\,
            I => \N__32283\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32280\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__32283\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__32280\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32266\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32266\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32266\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__32266\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32263\,
            I => \N__32260\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__32260\,
            I => \N__32257\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__32257\,
            I => \N__32254\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__32254\,
            I => \N__32251\
        );

    \I__5964\ : Odrv4
    port map (
            O => \N__32251\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32244\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__32247\,
            I => \N__32241\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32238\
        );

    \I__5960\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32234\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__32238\,
            I => \N__32231\
        );

    \I__5958\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32228\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__32234\,
            I => \N__32225\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__32231\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__32228\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__32225\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__32218\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \N__32212\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32208\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32205\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32202\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32199\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__32202\,
            I => \N__32196\
        );

    \I__5946\ : Span4Mux_h
    port map (
            O => \N__32199\,
            I => \N__32191\
        );

    \I__5945\ : Span4Mux_v
    port map (
            O => \N__32196\,
            I => \N__32191\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__32191\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32185\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32185\,
            I => \N__32180\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32177\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32174\
        );

    \I__5939\ : Span4Mux_h
    port map (
            O => \N__32180\,
            I => \N__32171\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32168\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__32174\,
            I => \N__32165\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__32171\,
            I => \N__32160\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__32168\,
            I => \N__32160\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__32165\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__32160\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__32155\,
            I => \N__32152\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32148\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__32151\,
            I => \N__32145\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32142\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32139\
        );

    \I__5927\ : Span4Mux_h
    port map (
            O => \N__32142\,
            I => \N__32133\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32139\,
            I => \N__32133\
        );

    \I__5925\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32130\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__32133\,
            I => \N__32126\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32123\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32120\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__32126\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__32123\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__32120\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32108\
        );

    \I__5917\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32105\
        );

    \I__5916\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32102\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__32108\,
            I => \N__32099\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32096\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32093\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__32099\,
            I => \N__32090\
        );

    \I__5911\ : Odrv12
    port map (
            O => \N__32096\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__32093\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__32090\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__32083\,
            I => \N__32080\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32077\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__32077\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__32074\,
            I => \N__32071\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32068\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__32068\,
            I => \N__32064\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32061\
        );

    \I__5901\ : Span4Mux_v
    port map (
            O => \N__32064\,
            I => \N__32056\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32056\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__32056\,
            I => \N__32053\
        );

    \I__5898\ : Span4Mux_h
    port map (
            O => \N__32053\,
            I => \N__32049\
        );

    \I__5897\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32046\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__32049\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__32046\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__32041\,
            I => \N__32038\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32034\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32037\,
            I => \N__32031\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__32034\,
            I => \N__32027\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__32031\,
            I => \N__32024\
        );

    \I__5889\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32020\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__32027\,
            I => \N__32017\
        );

    \I__5887\ : Span12Mux_v
    port map (
            O => \N__32024\,
            I => \N__32014\
        );

    \I__5886\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32011\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__32020\,
            I => \N__32008\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__32017\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5883\ : Odrv12
    port map (
            O => \N__32014\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__32011\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__32008\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__31999\,
            I => \N__31996\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31993\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__31993\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__31990\,
            I => \N__31986\
        );

    \I__5876\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31982\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31979\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31976\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31973\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31970\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31965\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__31973\,
            I => \N__31965\
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__31970\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__31965\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31953\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__31956\,
            I => \N__31949\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__31953\,
            I => \N__31946\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31943\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31939\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__31946\,
            I => \N__31934\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31934\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31931\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31939\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__31934\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31931\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__31924\,
            I => \N__31921\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31918\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31918\,
            I => \N__31915\
        );

    \I__5852\ : Span4Mux_h
    port map (
            O => \N__31915\,
            I => \N__31912\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__31912\,
            I => \N__31909\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__31909\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__31906\,
            I => \N__31903\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31900\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31897\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__31897\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31891\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__31888\,
            I => \N__31883\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31878\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31878\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__31883\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31878\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__31873\,
            I => \N__31869\
        );

    \I__5837\ : CascadeMux
    port map (
            O => \N__31872\,
            I => \N__31866\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31862\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31857\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31857\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31862\,
            I => \N__31854\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31857\,
            I => \N__31851\
        );

    \I__5831\ : Span12Mux_v
    port map (
            O => \N__31854\,
            I => \N__31847\
        );

    \I__5830\ : Span4Mux_h
    port map (
            O => \N__31851\,
            I => \N__31844\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31841\
        );

    \I__5828\ : Odrv12
    port map (
            O => \N__31847\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__31844\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31841\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__5825\ : CascadeMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31828\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31828\,
            I => \N__31825\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31822\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__31822\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31815\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31811\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31808\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__31814\,
            I => \N__31805\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31802\
        );

    \I__5815\ : Span4Mux_v
    port map (
            O => \N__31808\,
            I => \N__31799\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31796\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__31802\,
            I => \N__31793\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__31799\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31796\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__31793\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31783\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__31783\,
            I => \N__31779\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__31782\,
            I => \N__31775\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__31779\,
            I => \N__31772\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31769\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31766\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__31772\,
            I => \N__31761\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31761\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31757\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__31761\,
            I => \N__31754\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31751\
        );

    \I__5798\ : Odrv12
    port map (
            O => \N__31757\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__31754\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__31751\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31741\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__31735\,
            I => \N__31732\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__31732\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__31729\,
            I => \N__31726\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31723\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31719\
        );

    \I__5787\ : CascadeMux
    port map (
            O => \N__31722\,
            I => \N__31716\
        );

    \I__5786\ : Span4Mux_h
    port map (
            O => \N__31719\,
            I => \N__31712\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31709\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31706\
        );

    \I__5783\ : Span4Mux_v
    port map (
            O => \N__31712\,
            I => \N__31702\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31709\,
            I => \N__31699\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__31706\,
            I => \N__31696\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31705\,
            I => \N__31693\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__31702\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5778\ : Odrv12
    port map (
            O => \N__31699\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__31696\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__31693\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31679\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31676\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31673\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31670\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31667\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31664\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__31670\,
            I => \N__31661\
        );

    \I__5768\ : Odrv12
    port map (
            O => \N__31667\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__31664\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__31661\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__31654\,
            I => \N__31651\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31651\,
            I => \N__31648\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__31645\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__31642\,
            I => \N__31638\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31635\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31632\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__31635\,
            I => \N__31629\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31632\,
            I => \N__31623\
        );

    \I__5756\ : Span4Mux_v
    port map (
            O => \N__31629\,
            I => \N__31623\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31620\
        );

    \I__5754\ : Span4Mux_v
    port map (
            O => \N__31623\,
            I => \N__31616\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31613\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31610\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__31616\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__31613\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31610\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31595\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31592\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31589\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31586\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31592\,
            I => \N__31583\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31580\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__31586\,
            I => \N__31575\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__31583\,
            I => \N__31575\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__31580\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__31575\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31567\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31567\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__31564\,
            I => \N__31561\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31558\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__31558\,
            I => \N__31554\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31557\,
            I => \N__31551\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__31554\,
            I => \N__31547\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31544\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31541\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__31547\,
            I => \N__31538\
        );

    \I__5727\ : Span4Mux_v
    port map (
            O => \N__31544\,
            I => \N__31535\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__31541\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__31538\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__31535\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31524\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__31527\,
            I => \N__31520\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31524\,
            I => \N__31516\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31513\
        );

    \I__5719\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31508\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31508\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__31516\,
            I => \N__31503\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31503\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__31508\,
            I => \N__31500\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__31503\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__31500\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31489\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__31486\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__31483\,
            I => \N__31479\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__31482\,
            I => \N__31476\
        );

    \I__5706\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31472\
        );

    \I__5705\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31469\
        );

    \I__5704\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31466\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__31472\,
            I => \N__31461\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31461\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31458\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__31461\,
            I => \N__31454\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__31458\,
            I => \N__31451\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31448\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__31454\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__31451\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31448\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31438\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__31438\,
            I => \N__31434\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31431\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__31434\,
            I => \N__31425\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31431\,
            I => \N__31425\
        );

    \I__5689\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31422\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__31425\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__31422\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31414\
        );

    \I__5685\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31411\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31411\,
            I => \N__31408\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__31408\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__31405\,
            I => \N__31402\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31397\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31394\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31391\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31388\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__31394\,
            I => \N__31385\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__31391\,
            I => \N__31382\
        );

    \I__5675\ : Span4Mux_v
    port map (
            O => \N__31388\,
            I => \N__31379\
        );

    \I__5674\ : Span4Mux_v
    port map (
            O => \N__31385\,
            I => \N__31376\
        );

    \I__5673\ : Odrv12
    port map (
            O => \N__31382\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__31379\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__31376\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__31369\,
            I => \N__31366\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31362\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31359\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31355\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31352\
        );

    \I__5665\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31349\
        );

    \I__5664\ : Span4Mux_h
    port map (
            O => \N__31355\,
            I => \N__31345\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__31352\,
            I => \N__31340\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31340\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31337\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31334\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__31340\,
            I => \N__31331\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31328\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__31334\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__31331\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__31328\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31318\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__31318\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31312\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__31309\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31303\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31298\
        );

    \I__5647\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31295\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31292\
        );

    \I__5645\ : Span4Mux_v
    port map (
            O => \N__31298\,
            I => \N__31287\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__31295\,
            I => \N__31287\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31292\,
            I => \N__31283\
        );

    \I__5642\ : Span4Mux_h
    port map (
            O => \N__31287\,
            I => \N__31280\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31277\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__31283\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__31280\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__31277\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31265\
        );

    \I__5636\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31262\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__31268\,
            I => \N__31259\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31265\,
            I => \N__31256\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31253\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31250\
        );

    \I__5631\ : Span4Mux_v
    port map (
            O => \N__31256\,
            I => \N__31247\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__31253\,
            I => \N__31244\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__31250\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__31247\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__31244\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__31237\,
            I => \N__31234\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31231\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__31231\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__5623\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31223\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31217\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31217\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31214\
        );

    \I__5619\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31211\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31208\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__31214\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__31211\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__31208\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31196\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31193\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__31199\,
            I => \N__31190\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31187\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31184\
        );

    \I__5609\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31181\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__31187\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__31184\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31181\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__31174\,
            I => \N__31171\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31168\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31165\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__31165\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31158\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__31161\,
            I => \N__31155\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31158\,
            I => \N__31152\
        );

    \I__5598\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31149\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31146\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__31149\,
            I => \N__31143\
        );

    \I__5595\ : Span4Mux_v
    port map (
            O => \N__31146\,
            I => \N__31138\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__31143\,
            I => \N__31135\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31132\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31129\
        );

    \I__5591\ : Odrv4
    port map (
            O => \N__31138\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__31135\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__31132\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__31129\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__5587\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31116\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31113\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31110\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__31107\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__31110\,
            I => \N__31104\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__31107\,
            I => \N__31098\
        );

    \I__5581\ : Span4Mux_v
    port map (
            O => \N__31104\,
            I => \N__31098\
        );

    \I__5580\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31095\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__31098\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__31095\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__5577\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31087\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__31087\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__5575\ : InMux
    port map (
            O => \N__31084\,
            I => \N__31081\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31081\,
            I => \N__31076\
        );

    \I__5573\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31073\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31069\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__31076\,
            I => \N__31064\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31064\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31061\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N__31058\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__31064\,
            I => \N__31053\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__31061\,
            I => \N__31053\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__31058\,
            I => \N__31050\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__31053\,
            I => \N__31047\
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__31050\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__31047\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__5561\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31039\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__31039\,
            I => \N__31036\
        );

    \I__5559\ : Sp12to4
    port map (
            O => \N__31036\,
            I => \N__31033\
        );

    \I__5558\ : Odrv12
    port map (
            O => \N__31033\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__5557\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31026\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31023\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31020\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31017\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__31020\,
            I => \N__31014\
        );

    \I__5552\ : Span4Mux_s3_h
    port map (
            O => \N__31017\,
            I => \N__31011\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__31014\,
            I => \N__31008\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__31011\,
            I => \N__31005\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__31008\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__31005\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5547\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30997\,
            I => \N__30994\
        );

    \I__5545\ : Span4Mux_h
    port map (
            O => \N__30994\,
            I => \N__30991\
        );

    \I__5544\ : Odrv4
    port map (
            O => \N__30991\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__30988\,
            I => \N__30984\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__30987\,
            I => \N__30981\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30976\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30976\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30976\,
            I => \N__30973\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__30973\,
            I => \N__30968\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30963\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30963\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__30968\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__30963\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5533\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30952\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30952\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30952\,
            I => \N__30949\
        );

    \I__5530\ : Span4Mux_h
    port map (
            O => \N__30949\,
            I => \N__30945\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30942\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__30945\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__30942\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30934\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__30934\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__30931\,
            I => \N__30928\
        );

    \I__5523\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30925\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30922\
        );

    \I__5521\ : Span4Mux_h
    port map (
            O => \N__30922\,
            I => \N__30919\
        );

    \I__5520\ : Span4Mux_v
    port map (
            O => \N__30919\,
            I => \N__30916\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__30916\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__30913\,
            I => \N__30909\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30905\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30902\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30899\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__30905\,
            I => \N__30896\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__30902\,
            I => \N__30893\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30890\
        );

    \I__5511\ : Span4Mux_v
    port map (
            O => \N__30896\,
            I => \N__30885\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__30893\,
            I => \N__30885\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__30890\,
            I => \N__30882\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__30885\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__30882\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5506\ : CascadeMux
    port map (
            O => \N__30877\,
            I => \N__30874\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30871\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30871\,
            I => \N__30868\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__30868\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__30865\,
            I => \N__30861\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__30864\,
            I => \N__30858\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30855\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30851\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__30855\,
            I => \N__30848\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30845\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30851\,
            I => \N__30841\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__30848\,
            I => \N__30838\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30845\,
            I => \N__30835\
        );

    \I__5493\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30832\
        );

    \I__5492\ : Span4Mux_h
    port map (
            O => \N__30841\,
            I => \N__30829\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__30838\,
            I => \N__30826\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__30835\,
            I => \N__30821\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30821\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__30829\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__30826\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__30821\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30810\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30806\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30810\,
            I => \N__30803\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30800\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30806\,
            I => \N__30797\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__30803\,
            I => \N__30792\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30792\
        );

    \I__5478\ : Span4Mux_v
    port map (
            O => \N__30797\,
            I => \N__30789\
        );

    \I__5477\ : Span4Mux_v
    port map (
            O => \N__30792\,
            I => \N__30786\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__30789\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__30786\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__30781\,
            I => \N__30778\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30775\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30775\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__30772\,
            I => \N__30769\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30765\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30762\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30758\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30755\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30752\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__30758\,
            I => \N__30748\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30743\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30752\,
            I => \N__30743\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30751\,
            I => \N__30740\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__30748\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__30743\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30740\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30733\,
            I => \N__30730\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30730\,
            I => \N__30725\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30720\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30720\
        );

    \I__5454\ : Span4Mux_v
    port map (
            O => \N__30725\,
            I => \N__30717\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30720\,
            I => \N__30714\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__30717\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__30714\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30709\,
            I => \N__30706\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30703\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30703\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__30700\,
            I => \N__30697\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30691\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30691\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30691\,
            I => \N__30688\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30685\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__30685\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30679\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__30679\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__30670\,
            I => \N__30665\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30660\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30660\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__30665\,
            I => \N__30654\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30660\,
            I => \N__30654\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30651\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__30654\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30651\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30643\,
            I => \N__30640\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__30640\,
            I => \N__30636\
        );

    \I__5426\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30633\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__30636\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30633\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30622\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30622\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30622\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30614\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30608\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30608\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30614\,
            I => \N__30605\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30602\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30599\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__30605\,
            I => \N__30596\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30593\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__30599\,
            I => \N__30590\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__30596\,
            I => \N__30585\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__30593\,
            I => \N__30585\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__30590\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__30585\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30577\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__30577\,
            I => \N__30574\
        );

    \I__5405\ : Span4Mux_v
    port map (
            O => \N__30574\,
            I => \N__30570\
        );

    \I__5404\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30567\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__30570\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__30567\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__5401\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30543\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30543\
        );

    \I__5399\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30538\
        );

    \I__5398\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30538\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__30558\,
            I => \N__30531\
        );

    \I__5396\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30523\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30516\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30516\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30516\
        );

    \I__5392\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30505\
        );

    \I__5391\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30505\
        );

    \I__5390\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30505\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30505\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30505\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__30548\,
            I => \N__30494\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30487\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__30538\,
            I => \N__30484\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30467\
        );

    \I__5383\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30467\
        );

    \I__5382\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30467\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30467\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30467\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30467\
        );

    \I__5378\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30467\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30467\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30462\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30462\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30455\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30455\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__30505\,
            I => \N__30455\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30442\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30442\
        );

    \I__5369\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30442\
        );

    \I__5368\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30442\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30442\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30442\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30416\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30409\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30409\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30409\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30402\
        );

    \I__5360\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30402\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30402\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__30487\,
            I => \N__30389\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__30484\,
            I => \N__30389\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__30467\,
            I => \N__30389\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30389\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__30455\,
            I => \N__30389\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__30442\,
            I => \N__30389\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30378\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30378\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30378\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30378\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30378\
        );

    \I__5347\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30369\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30369\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30369\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30369\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30365\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30358\
        );

    \I__5341\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30358\
        );

    \I__5340\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30358\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30347\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30347\
        );

    \I__5337\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30347\
        );

    \I__5336\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30347\
        );

    \I__5335\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30343\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30336\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30336\
        );

    \I__5332\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30336\
        );

    \I__5331\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30331\
        );

    \I__5330\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30331\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__30416\,
            I => \N__30306\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__30409\,
            I => \N__30306\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30306\
        );

    \I__5326\ : Span4Mux_h
    port map (
            O => \N__30389\,
            I => \N__30306\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__30378\,
            I => \N__30306\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30306\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30299\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30296\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__30358\,
            I => \N__30293\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30288\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30288\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30285\
        );

    \I__5317\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30282\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N__30275\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__30336\,
            I => \N__30275\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__30331\,
            I => \N__30275\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30330\,
            I => \N__30270\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30270\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30267\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30260\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30260\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30325\,
            I => \N__30260\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30255\
        );

    \I__5306\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30255\
        );

    \I__5305\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30248\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30248\
        );

    \I__5303\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30248\
        );

    \I__5302\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30238\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__30306\,
            I => \N__30235\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30228\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30228\
        );

    \I__5298\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30228\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30222\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__30299\,
            I => \N__30210\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__30296\,
            I => \N__30210\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__30293\,
            I => \N__30210\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30288\,
            I => \N__30210\
        );

    \I__5292\ : Span4Mux_v
    port map (
            O => \N__30285\,
            I => \N__30205\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__30282\,
            I => \N__30205\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__30275\,
            I => \N__30198\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__30270\,
            I => \N__30198\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30198\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30191\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__30255\,
            I => \N__30191\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__30248\,
            I => \N__30191\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30188\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30183\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30183\
        );

    \I__5281\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30180\
        );

    \I__5280\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30177\
        );

    \I__5279\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30172\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30172\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__30238\,
            I => \N__30165\
        );

    \I__5276\ : Sp12to4
    port map (
            O => \N__30235\,
            I => \N__30165\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__30228\,
            I => \N__30165\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30160\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30160\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30225\,
            I => \N__30157\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30222\,
            I => \N__30154\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30147\
        );

    \I__5269\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30147\
        );

    \I__5268\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30147\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__30210\,
            I => \N__30142\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__30205\,
            I => \N__30142\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__30198\,
            I => \N__30139\
        );

    \I__5264\ : Span12Mux_v
    port map (
            O => \N__30191\,
            I => \N__30136\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30123\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__30183\,
            I => \N__30123\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__30180\,
            I => \N__30123\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__30177\,
            I => \N__30123\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30123\
        );

    \I__5258\ : Span12Mux_h
    port map (
            O => \N__30165\,
            I => \N__30123\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30160\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__30157\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__30154\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__30147\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__30142\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__30139\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__30136\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__30123\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__5249\ : CEMux
    port map (
            O => \N__30106\,
            I => \N__30073\
        );

    \I__5248\ : CEMux
    port map (
            O => \N__30105\,
            I => \N__30073\
        );

    \I__5247\ : CEMux
    port map (
            O => \N__30104\,
            I => \N__30073\
        );

    \I__5246\ : CEMux
    port map (
            O => \N__30103\,
            I => \N__30073\
        );

    \I__5245\ : CEMux
    port map (
            O => \N__30102\,
            I => \N__30073\
        );

    \I__5244\ : CEMux
    port map (
            O => \N__30101\,
            I => \N__30073\
        );

    \I__5243\ : CEMux
    port map (
            O => \N__30100\,
            I => \N__30073\
        );

    \I__5242\ : CEMux
    port map (
            O => \N__30099\,
            I => \N__30073\
        );

    \I__5241\ : CEMux
    port map (
            O => \N__30098\,
            I => \N__30073\
        );

    \I__5240\ : CEMux
    port map (
            O => \N__30097\,
            I => \N__30073\
        );

    \I__5239\ : CEMux
    port map (
            O => \N__30096\,
            I => \N__30073\
        );

    \I__5238\ : GlobalMux
    port map (
            O => \N__30073\,
            I => \N__30070\
        );

    \I__5237\ : gio2CtrlBuf
    port map (
            O => \N__30070\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30064\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__30064\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__30061\,
            I => \N__30058\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30052\
        );

    \I__5232\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30052\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__30052\,
            I => \N__30049\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__30046\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__5228\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30037\
        );

    \I__5227\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30037\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__30037\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30028\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__30028\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30022\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__30022\,
            I => \N__30018\
        );

    \I__5220\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30015\
        );

    \I__5219\ : Span4Mux_h
    port map (
            O => \N__30018\,
            I => \N__30010\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__30010\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__30010\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__30007\,
            I => \N__30003\
        );

    \I__5215\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30000\
        );

    \I__5214\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29997\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__30000\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__29997\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__29986\,
            I => \N__29983\
        );

    \I__5208\ : Odrv4
    port map (
            O => \N__29983\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__5207\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29976\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29973\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29976\,
            I => \N__29970\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29973\,
            I => \N__29967\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__29970\,
            I => \N__29964\
        );

    \I__5202\ : Span12Mux_v
    port map (
            O => \N__29967\,
            I => \N__29961\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__29964\,
            I => \N__29958\
        );

    \I__5200\ : Odrv12
    port map (
            O => \N__29961\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__29958\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29950\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29950\,
            I => \N__29946\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29943\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__29946\,
            I => \N__29940\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29937\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__29940\,
            I => \N__29934\
        );

    \I__5192\ : Span12Mux_s7_h
    port map (
            O => \N__29937\,
            I => \N__29931\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__29934\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5190\ : Odrv12
    port map (
            O => \N__29931\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29922\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29919\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29916\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29919\,
            I => \N__29913\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__29916\,
            I => \N__29910\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__29913\,
            I => \N__29907\
        );

    \I__5183\ : Sp12to4
    port map (
            O => \N__29910\,
            I => \N__29904\
        );

    \I__5182\ : Sp12to4
    port map (
            O => \N__29907\,
            I => \N__29899\
        );

    \I__5181\ : Span12Mux_v
    port map (
            O => \N__29904\,
            I => \N__29899\
        );

    \I__5180\ : Odrv12
    port map (
            O => \N__29899\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__29893\,
            I => \N__29890\
        );

    \I__5177\ : Odrv12
    port map (
            O => \N__29890\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29881\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29878\
        );

    \I__5173\ : Odrv12
    port map (
            O => \N__29878\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29872\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__29872\,
            I => \N__29869\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__29869\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__29866\,
            I => \N__29863\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29860\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__29860\,
            I => \N__29857\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__29857\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29851\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29851\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__29848\,
            I => \N__29845\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29842\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29842\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29836\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29836\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29833\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__29830\,
            I => \N__29827\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29824\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__29824\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__29821\,
            I => \N__29818\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29815\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29815\,
            I => \N__29812\
        );

    \I__5151\ : Odrv12
    port map (
            O => \N__29812\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29806\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29806\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29797\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__29794\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29788\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29788\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29782\,
            I => \N__29779\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__29779\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__29776\,
            I => \N__29773\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29770\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29770\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29764\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29764\,
            I => \N__29761\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__29761\,
            I => \N__29758\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__29758\,
            I => \N__29755\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__29755\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__29752\,
            I => \N__29749\
        );

    \I__5130\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29746\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29740\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29740\,
            I => \N__29737\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__29737\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29728\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__29728\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__5122\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29719\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__29719\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__29716\,
            I => \N__29713\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29710\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29710\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29704\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29695\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__29695\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29689\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29689\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29680\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__29677\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__5105\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29671\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__29671\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__29668\,
            I => \N__29665\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__29662\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29656\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29656\,
            I => \N__29653\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__29653\,
            I => \N__29650\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__29650\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__29647\,
            I => \N__29644\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__29641\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29635\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29632\
        );

    \I__5091\ : Odrv12
    port map (
            O => \N__29632\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__29629\,
            I => \N__29626\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29623\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__29623\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29617\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29617\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__29614\,
            I => \N__29611\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29608\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29605\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__29605\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__29602\,
            I => \N__29599\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29599\,
            I => \N__29596\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__29596\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29590\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__29581\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29575\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__29572\,
            I => \N__29569\
        );

    \I__5070\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29566\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__29566\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29560\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29560\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__29554\,
            I => \N__29551\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__29551\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__5062\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29542\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__29542\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29534\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29531\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29528\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29534\,
            I => \N__29523\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29531\,
            I => \N__29523\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29528\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__29523\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29514\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29511\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__29514\,
            I => \N__29508\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__29511\,
            I => \N__29504\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__29508\,
            I => \N__29501\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29498\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__29504\,
            I => \N__29495\
        );

    \I__5046\ : Sp12to4
    port map (
            O => \N__29501\,
            I => \N__29489\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29489\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__29495\,
            I => \N__29486\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29483\
        );

    \I__5042\ : Odrv12
    port map (
            O => \N__29489\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__29486\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__29483\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__29476\,
            I => \N__29472\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29467\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29467\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29467\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__5035\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29459\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29463\,
            I => \N__29454\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29454\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29451\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29448\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__29448\,
            I => \N__29442\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29439\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__29442\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29439\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5025\ : InMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__29431\,
            I => \N__29427\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29424\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__29427\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__29424\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5020\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29413\
        );

    \I__5019\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29413\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29413\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29407\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29407\,
            I => \N__29403\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29400\
        );

    \I__5014\ : Odrv4
    port map (
            O => \N__29403\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29400\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__5012\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29390\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29385\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29385\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29379\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29379\
        );

    \I__5007\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29376\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__29379\,
            I => \N__29371\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__29376\,
            I => \N__29371\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__29368\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5002\ : CascadeMux
    port map (
            O => \N__29365\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29357\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29352\
        );

    \I__4999\ : InMux
    port map (
            O => \N__29360\,
            I => \N__29352\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29357\,
            I => \N__29346\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__29352\,
            I => \N__29346\
        );

    \I__4996\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29343\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__29346\,
            I => \N__29338\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__29343\,
            I => \N__29338\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__29338\,
            I => \N__29335\
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__29335\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29328\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29325\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29328\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__29325\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__29320\,
            I => \N__29317\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29314\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29314\,
            I => \N__29311\
        );

    \I__4984\ : Odrv12
    port map (
            O => \N__29311\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__4983\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29305\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__29305\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__29302\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29296\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29296\,
            I => \N__29293\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__29293\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__29290\,
            I => \N__29287\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29284\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__29284\,
            I => \N__29281\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__29281\,
            I => \N__29278\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__29278\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__4972\ : CEMux
    port map (
            O => \N__29275\,
            I => \N__29271\
        );

    \I__4971\ : CEMux
    port map (
            O => \N__29274\,
            I => \N__29268\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29260\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29260\
        );

    \I__4968\ : CEMux
    port map (
            O => \N__29267\,
            I => \N__29257\
        );

    \I__4967\ : CEMux
    port map (
            O => \N__29266\,
            I => \N__29249\
        );

    \I__4966\ : CEMux
    port map (
            O => \N__29265\,
            I => \N__29243\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__29260\,
            I => \N__29230\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29230\
        );

    \I__4963\ : CEMux
    port map (
            O => \N__29256\,
            I => \N__29227\
        );

    \I__4962\ : CEMux
    port map (
            O => \N__29255\,
            I => \N__29220\
        );

    \I__4961\ : CEMux
    port map (
            O => \N__29254\,
            I => \N__29216\
        );

    \I__4960\ : CEMux
    port map (
            O => \N__29253\,
            I => \N__29212\
        );

    \I__4959\ : CEMux
    port map (
            O => \N__29252\,
            I => \N__29209\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__29249\,
            I => \N__29206\
        );

    \I__4957\ : CEMux
    port map (
            O => \N__29248\,
            I => \N__29203\
        );

    \I__4956\ : CEMux
    port map (
            O => \N__29247\,
            I => \N__29200\
        );

    \I__4955\ : CEMux
    port map (
            O => \N__29246\,
            I => \N__29197\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29183\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29174\
        );

    \I__4952\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29174\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29174\
        );

    \I__4950\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29174\
        );

    \I__4949\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29167\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29167\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29167\
        );

    \I__4946\ : CEMux
    port map (
            O => \N__29235\,
            I => \N__29164\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__29230\,
            I => \N__29159\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29159\
        );

    \I__4943\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29150\
        );

    \I__4942\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29150\
        );

    \I__4941\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29150\
        );

    \I__4940\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29150\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29146\
        );

    \I__4938\ : CEMux
    port map (
            O => \N__29219\,
            I => \N__29143\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29216\,
            I => \N__29140\
        );

    \I__4936\ : CEMux
    port map (
            O => \N__29215\,
            I => \N__29137\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__29212\,
            I => \N__29132\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29132\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__29206\,
            I => \N__29125\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29203\,
            I => \N__29125\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29125\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29114\
        );

    \I__4929\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29105\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29105\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29105\
        );

    \I__4926\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29105\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29098\
        );

    \I__4924\ : InMux
    port map (
            O => \N__29191\,
            I => \N__29098\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29098\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29089\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29089\
        );

    \I__4920\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29089\
        );

    \I__4919\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29089\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__29183\,
            I => \N__29082\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29082\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__29167\,
            I => \N__29082\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__29164\,
            I => \N__29077\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__29159\,
            I => \N__29077\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29074\
        );

    \I__4912\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29071\
        );

    \I__4911\ : Span4Mux_h
    port map (
            O => \N__29146\,
            I => \N__29068\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__29143\,
            I => \N__29063\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__29140\,
            I => \N__29063\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__29137\,
            I => \N__29058\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__29132\,
            I => \N__29058\
        );

    \I__4906\ : Span4Mux_v
    port map (
            O => \N__29125\,
            I => \N__29055\
        );

    \I__4905\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29046\
        );

    \I__4904\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29046\
        );

    \I__4903\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29046\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29046\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29037\
        );

    \I__4900\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29037\
        );

    \I__4899\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29037\
        );

    \I__4898\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29037\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__29114\,
            I => \N__29034\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29031\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29020\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29020\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__29082\,
            I => \N__29020\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__29077\,
            I => \N__29020\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__29074\,
            I => \N__29020\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__29071\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__29068\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__29063\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__29058\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__29055\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__29046\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__29037\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__29034\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__29031\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__29020\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28996\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__28996\,
            I => \N__28991\
        );

    \I__4878\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28988\
        );

    \I__4877\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28985\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__28991\,
            I => \N__28982\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28979\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28976\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__28982\,
            I => \N__28970\
        );

    \I__4872\ : Span4Mux_h
    port map (
            O => \N__28979\,
            I => \N__28970\
        );

    \I__4871\ : Span12Mux_h
    port map (
            O => \N__28976\,
            I => \N__28967\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28964\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__28970\,
            I => \N__28961\
        );

    \I__4868\ : Span12Mux_v
    port map (
            O => \N__28967\,
            I => \N__28958\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__28964\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__28961\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4865\ : Odrv12
    port map (
            O => \N__28958\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__4864\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28948\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28942\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28935\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28935\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28935\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__28942\,
            I => \N__28930\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28935\,
            I => \N__28930\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__28930\,
            I => \N__28927\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__28927\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28921\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__28921\,
            I => \N__28917\
        );

    \I__4853\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28914\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__28917\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28914\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28904\
        );

    \I__4849\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28899\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28899\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28893\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28893\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28890\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28885\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__28885\,
            I => \N__28882\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__28882\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28875\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28872\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__28875\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28872\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4836\ : InMux
    port map (
            O => \N__28867\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28860\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__28863\,
            I => \N__28857\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28860\,
            I => \N__28853\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28850\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28847\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__28853\,
            I => \N__28844\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28850\,
            I => \N__28841\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28838\
        );

    \I__4827\ : Span4Mux_v
    port map (
            O => \N__28844\,
            I => \N__28832\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__28841\,
            I => \N__28832\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__28838\,
            I => \N__28829\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28826\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__28832\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__28829\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28826\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__28819\,
            I => \N__28815\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28812\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28809\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28812\,
            I => \N__28805\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28802\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28799\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__28805\,
            I => \N__28796\
        );

    \I__4813\ : Odrv12
    port map (
            O => \N__28802\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__28799\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__28796\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28783\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28780\
        );

    \I__4807\ : Odrv12
    port map (
            O => \N__28780\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28765\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28762\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28757\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28757\
        );

    \I__4800\ : Span4Mux_v
    port map (
            O => \N__28765\,
            I => \N__28754\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28762\,
            I => \N__28751\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28748\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__28754\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__28751\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__28748\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__28740\,
            I => \N__28734\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28737\,
            I => \N__28730\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28727\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28724\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__28730\,
            I => \N__28721\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28727\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28724\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__28721\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__28714\,
            I => \N__28711\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28708\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28708\,
            I => \N__28705\
        );

    \I__4782\ : Odrv12
    port map (
            O => \N__28705\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__4781\ : IoInMux
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__28699\,
            I => \N__28696\
        );

    \I__4779\ : IoSpan4Mux
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__4778\ : Span4Mux_s0_v
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__28690\,
            I => s3_phy_c
        );

    \I__4776\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__4774\ : Glb2LocalMux
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__4773\ : GlobalMux
    port map (
            O => \N__28678\,
            I => clk_12mhz
        );

    \I__4772\ : IoInMux
    port map (
            O => \N__28675\,
            I => \N__28672\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28672\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28664\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28661\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28658\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28664\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28661\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__28658\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28647\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28643\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28647\,
            I => \N__28640\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28637\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28643\,
            I => \N__28633\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__28640\,
            I => \N__28628\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28628\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__28636\,
            I => \N__28625\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__28633\,
            I => \N__28622\
        );

    \I__4755\ : Span4Mux_h
    port map (
            O => \N__28628\,
            I => \N__28619\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28616\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__28622\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__28619\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28616\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28606\,
            I => \N__28600\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28595\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28595\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28592\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__28600\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28595\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__28592\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__28585\,
            I => \N__28581\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__28584\,
            I => \N__28578\
        );

    \I__4740\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28572\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28569\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28562\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28562\
        );

    \I__4736\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28562\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__28572\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28569\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__28562\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28551\
        );

    \I__4731\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28548\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28542\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28542\
        );

    \I__4728\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28539\
        );

    \I__4727\ : Span4Mux_h
    port map (
            O => \N__28542\,
            I => \N__28536\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__28536\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__4724\ : Odrv12
    port map (
            O => \N__28533\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28525\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__28525\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28519\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28515\
        );

    \I__4719\ : InMux
    port map (
            O => \N__28518\,
            I => \N__28512\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28506\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__28512\,
            I => \N__28506\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28503\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__28506\,
            I => \N__28500\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28503\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__28500\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28495\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__28489\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28486\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__28480\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28477\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28471\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__4703\ : InMux
    port map (
            O => \N__28468\,
            I => \bfn_11_25_0_\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28462\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28456\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28456\,
            I => \N__28452\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__28455\,
            I => \N__28449\
        );

    \I__4697\ : Span4Mux_h
    port map (
            O => \N__28452\,
            I => \N__28446\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28442\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__28446\,
            I => \N__28439\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28436\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28442\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__28439\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__28436\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28429\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__4689\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28420\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__28420\,
            I => \N__28417\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__28417\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28414\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28411\,
            I => \N__28408\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__28408\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__4682\ : InMux
    port map (
            O => \N__28405\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__4681\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28399\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__28399\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28396\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28390\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__28390\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__28387\,
            I => \N__28384\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28377\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28377\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28374\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28377\,
            I => \N__28371\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28368\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__28371\,
            I => \N__28365\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__28368\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__28365\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__4667\ : InMux
    port map (
            O => \N__28360\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__4666\ : InMux
    port map (
            O => \N__28357\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28354\,
            I => \N__28351\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28351\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__4663\ : InMux
    port map (
            O => \N__28348\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__4662\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28342\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__28342\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28339\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__4659\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__4657\ : Odrv12
    port map (
            O => \N__28330\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28327\,
            I => \bfn_11_24_0_\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28321\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28318\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28312\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__28312\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28309\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28303\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__28303\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28296\
        );

    \I__4646\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28293\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28285\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__28290\,
            I => \N__28285\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__28285\,
            I => \N__28281\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28278\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__28281\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28278\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4638\ : InMux
    port map (
            O => \N__28273\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__4637\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28267\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28267\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28264\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__4634\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28258\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__28258\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__28255\,
            I => \N__28251\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__28254\,
            I => \N__28248\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28245\
        );

    \I__4629\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28242\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28238\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__28242\,
            I => \N__28235\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28232\
        );

    \I__4625\ : Span4Mux_h
    port map (
            O => \N__28238\,
            I => \N__28227\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__28235\,
            I => \N__28227\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__28232\,
            I => \N__28224\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__28227\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__4621\ : Odrv12
    port map (
            O => \N__28224\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__4620\ : InMux
    port map (
            O => \N__28219\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28213\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__4617\ : InMux
    port map (
            O => \N__28210\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28201\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__28201\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__4613\ : InMux
    port map (
            O => \N__28198\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28189\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__28189\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__4609\ : InMux
    port map (
            O => \N__28186\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28180\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28177\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__28177\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28174\,
            I => \bfn_11_23_0_\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28168\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__28168\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__4602\ : InMux
    port map (
            O => \N__28165\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__4601\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28159\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__28159\,
            I => \N__28156\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__28153\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28150\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__4596\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28144\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__28144\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28141\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28135\,
            I => \N__28132\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__28132\,
            I => \N__28129\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__28129\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__4589\ : InMux
    port map (
            O => \N__28126\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__4588\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28120\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__28120\,
            I => \N__28117\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__28117\,
            I => \N__28114\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__28114\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28111\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28102\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__28102\,
            I => \N__28099\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__28099\,
            I => \N__28096\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__28096\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__4578\ : InMux
    port map (
            O => \N__28093\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__4577\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28087\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__28087\,
            I => \N__28084\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__28084\,
            I => \N__28081\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__28081\,
            I => \N__28078\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__28078\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__4572\ : InMux
    port map (
            O => \N__28075\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28072\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28066\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28063\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__28063\,
            I => \N__28060\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__28060\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__4566\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28054\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__28054\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__4564\ : InMux
    port map (
            O => \N__28051\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__4563\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__28045\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28042\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28036\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__28036\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__4558\ : InMux
    port map (
            O => \N__28033\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__4557\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28027\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__28027\,
            I => \N__28024\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__4554\ : Sp12to4
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__4553\ : Odrv12
    port map (
            O => \N__28018\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__4552\ : InMux
    port map (
            O => \N__28015\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__4550\ : InMux
    port map (
            O => \N__28009\,
            I => \N__28006\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__28006\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28003\,
            I => \N__28000\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__27994\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27991\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27985\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27982\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__27982\,
            I => \N__27979\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__27979\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27976\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__27973\,
            I => \N__27970\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27967\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__27967\,
            I => \N__27964\
        );

    \I__4535\ : Span12Mux_v
    port map (
            O => \N__27964\,
            I => \N__27961\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__27961\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__27955\,
            I => \N__27952\
        );

    \I__4531\ : Span4Mux_v
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__27949\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27946\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27940\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__4526\ : Span12Mux_s11_h
    port map (
            O => \N__27937\,
            I => \N__27934\
        );

    \I__4525\ : Odrv12
    port map (
            O => \N__27934\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27931\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27925\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__27925\,
            I => \N__27922\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__27922\,
            I => \N__27919\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__27919\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27916\,
            I => \bfn_11_21_0_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27910\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27907\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__27907\,
            I => \N__27904\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__27904\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27901\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__27898\,
            I => \N__27895\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27892\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27889\
        );

    \I__4510\ : Span4Mux_h
    port map (
            O => \N__27889\,
            I => \N__27886\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__27886\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27880\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27877\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__27877\,
            I => \N__27874\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__27874\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27871\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__4501\ : Span4Mux_v
    port map (
            O => \N__27862\,
            I => \N__27859\
        );

    \I__4500\ : Span4Mux_v
    port map (
            O => \N__27859\,
            I => \N__27856\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__27856\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27853\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__27847\,
            I => \N__27844\
        );

    \I__4495\ : Span4Mux_h
    port map (
            O => \N__27844\,
            I => \N__27841\
        );

    \I__4494\ : Sp12to4
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__27838\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27835\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27829\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27823\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27823\,
            I => \N__27820\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__27820\,
            I => \N__27817\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__27817\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27814\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__4482\ : Span12Mux_v
    port map (
            O => \N__27805\,
            I => \N__27802\
        );

    \I__4481\ : Odrv12
    port map (
            O => \N__27802\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27799\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27793\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27790\
        );

    \I__4477\ : Span4Mux_h
    port map (
            O => \N__27790\,
            I => \N__27787\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__27784\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27781\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27775\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27772\
        );

    \I__4471\ : Span4Mux_v
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__4470\ : Span4Mux_v
    port map (
            O => \N__27769\,
            I => \N__27766\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__27766\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27763\,
            I => \bfn_11_20_0_\
        );

    \I__4467\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27757\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27754\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__27754\,
            I => \N__27751\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__27751\,
            I => \N__27748\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__27745\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__4461\ : InMux
    port map (
            O => \N__27742\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27736\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__27736\,
            I => \N__27733\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__27733\,
            I => \N__27730\
        );

    \I__4457\ : Span4Mux_v
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__27727\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27724\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__4454\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27718\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27718\,
            I => \N__27715\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__27712\,
            I => \N__27709\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__27709\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27706\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27700\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27697\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__27694\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27691\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__27685\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27679\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__27679\,
            I => \N__27676\
        );

    \I__4439\ : Span4Mux_h
    port map (
            O => \N__27676\,
            I => \N__27673\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__27673\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27670\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__27664\,
            I => \N__27661\
        );

    \I__4434\ : Span12Mux_v
    port map (
            O => \N__27661\,
            I => \N__27658\
        );

    \I__4433\ : Odrv12
    port map (
            O => \N__27658\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27655\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27649\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27649\,
            I => \N__27646\
        );

    \I__4429\ : Span4Mux_h
    port map (
            O => \N__27646\,
            I => \N__27643\
        );

    \I__4428\ : Span4Mux_v
    port map (
            O => \N__27643\,
            I => \N__27640\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__27640\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27637\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27631\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27631\,
            I => \N__27628\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__27628\,
            I => \N__27625\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__27625\,
            I => \N__27622\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__27622\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27619\,
            I => \bfn_11_19_0_\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27613\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27613\,
            I => \N__27610\
        );

    \I__4417\ : Span4Mux_h
    port map (
            O => \N__27610\,
            I => \N__27607\
        );

    \I__4416\ : Sp12to4
    port map (
            O => \N__27607\,
            I => \N__27604\
        );

    \I__4415\ : Span12Mux_v
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__27601\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27598\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27592\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27589\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__27589\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27586\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27583\,
            I => \N__27580\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__27580\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__4406\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27574\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__4404\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27568\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27568\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__27565\,
            I => \N__27562\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27559\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27559\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27553\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27553\,
            I => \N__27550\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__27550\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__27547\,
            I => \N__27544\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27541\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27541\,
            I => \N__27538\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__27538\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__27535\,
            I => \N__27532\
        );

    \I__4391\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27529\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27526\
        );

    \I__4389\ : Span4Mux_h
    port map (
            O => \N__27526\,
            I => \N__27522\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27519\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__27522\,
            I => \N__27514\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__27519\,
            I => \N__27514\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__27514\,
            I => \N__27511\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__27511\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__27508\,
            I => \N__27505\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27502\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27502\,
            I => \N__27498\
        );

    \I__4380\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27495\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__27498\,
            I => \N__27492\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27495\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__27492\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__27487\,
            I => \N__27484\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27481\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27481\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__4373\ : InMux
    port map (
            O => \N__27478\,
            I => \N__27475\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__27475\,
            I => \N__27470\
        );

    \I__4371\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27466\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27463\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__27470\,
            I => \N__27460\
        );

    \I__4368\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27457\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__27466\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27463\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__27460\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27457\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__27448\,
            I => \N__27445\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27442\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27439\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__27439\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27430\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27430\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__27427\,
            I => \N__27424\
        );

    \I__4355\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27421\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__27418\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__27415\,
            I => \N__27412\
        );

    \I__4351\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27408\
        );

    \I__4350\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27404\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27401\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__27407\,
            I => \N__27398\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27395\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__27401\,
            I => \N__27392\
        );

    \I__4345\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27389\
        );

    \I__4344\ : Span4Mux_v
    port map (
            O => \N__27395\,
            I => \N__27386\
        );

    \I__4343\ : Span4Mux_v
    port map (
            O => \N__27392\,
            I => \N__27382\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27389\,
            I => \N__27377\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__27386\,
            I => \N__27377\
        );

    \I__4340\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27374\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__27382\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__27377\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__27374\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__27367\,
            I => \N__27364\
        );

    \I__4335\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__27361\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27352\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27352\,
            I => \N__27349\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__27349\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27343\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__27343\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27337\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27334\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__27334\,
            I => \N__27331\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__27331\,
            I => \N__27326\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27323\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27319\
        );

    \I__4321\ : Span4Mux_h
    port map (
            O => \N__27326\,
            I => \N__27314\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27314\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27311\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27319\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__4317\ : Odrv4
    port map (
            O => \N__27314\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27311\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__27304\,
            I => \N__27301\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27298\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__27298\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__27295\,
            I => \N__27292\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27289\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27289\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27283\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27283\,
            I => \N__27278\
        );

    \I__4307\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27273\
        );

    \I__4306\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27273\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__27278\,
            I => \N__27268\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__27273\,
            I => \N__27268\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__27268\,
            I => \N__27264\
        );

    \I__4302\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27261\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__27264\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__27261\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__27253\,
            I => \N__27249\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27246\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__27249\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__27246\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4294\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27235\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27235\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27235\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27227\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27224\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27221\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27227\,
            I => \N__27218\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__27224\,
            I => \N__27215\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__27221\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4285\ : Odrv12
    port map (
            O => \N__27218\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__27215\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4283\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27203\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27200\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27197\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27194\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__27200\,
            I => \N__27191\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27197\,
            I => \N__27188\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__27194\,
            I => \N__27184\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__27191\,
            I => \N__27179\
        );

    \I__4275\ : Span4Mux_h
    port map (
            O => \N__27188\,
            I => \N__27179\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27176\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__27184\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__27179\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27176\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__27169\,
            I => \N__27166\
        );

    \I__4269\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27160\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27165\,
            I => \N__27160\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__27160\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__4265\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27148\
        );

    \I__4264\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27145\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27140\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27140\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27135\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27145\,
            I => \N__27135\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27132\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__27135\,
            I => \N__27129\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__27132\,
            I => \N__27126\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__27129\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__27126\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4254\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27118\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__27118\,
            I => \N__27113\
        );

    \I__4252\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27110\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27107\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__27113\,
            I => \N__27104\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__27110\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27107\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__27104\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27091\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27088\
        );

    \I__4243\ : Odrv12
    port map (
            O => \N__27088\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__4242\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27082\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27077\
        );

    \I__4240\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27074\
        );

    \I__4239\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27071\
        );

    \I__4238\ : Span4Mux_h
    port map (
            O => \N__27077\,
            I => \N__27068\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27065\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__27071\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__27068\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4234\ : Odrv12
    port map (
            O => \N__27065\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27054\
        );

    \I__4232\ : InMux
    port map (
            O => \N__27057\,
            I => \N__27050\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__27054\,
            I => \N__27047\
        );

    \I__4230\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27044\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27041\
        );

    \I__4228\ : Span4Mux_v
    port map (
            O => \N__27047\,
            I => \N__27037\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27044\,
            I => \N__27034\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__27041\,
            I => \N__27031\
        );

    \I__4225\ : InMux
    port map (
            O => \N__27040\,
            I => \N__27028\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__27037\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__27034\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__27031\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__27028\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__27019\,
            I => \N__27016\
        );

    \I__4219\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27010\
        );

    \I__4218\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27010\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27010\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__4216\ : InMux
    port map (
            O => \N__27007\,
            I => \N__27003\
        );

    \I__4215\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26998\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26995\
        );

    \I__4213\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26990\
        );

    \I__4212\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26990\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26987\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__26995\,
            I => \N__26982\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26982\
        );

    \I__4208\ : Span4Mux_h
    port map (
            O => \N__26987\,
            I => \N__26979\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__26982\,
            I => \N__26976\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__26979\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__26976\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26968\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26968\,
            I => \N__26964\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26960\
        );

    \I__4201\ : Span12Mux_h
    port map (
            O => \N__26964\,
            I => \N__26957\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26954\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__26960\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4198\ : Odrv12
    port map (
            O => \N__26957\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26954\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4196\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__26944\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26938\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26935\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__26935\,
            I => \N__26931\
        );

    \I__4191\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26927\
        );

    \I__4190\ : Span4Mux_v
    port map (
            O => \N__26931\,
            I => \N__26924\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26921\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__26927\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__26924\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__26921\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26908\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26905\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26902\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26899\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26896\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__26905\,
            I => \N__26893\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26902\,
            I => \N__26890\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26887\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__26896\,
            I => \N__26880\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__26893\,
            I => \N__26880\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__26890\,
            I => \N__26880\
        );

    \I__4174\ : Odrv12
    port map (
            O => \N__26887\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__26880\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__4172\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26869\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26869\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26869\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26862\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__26865\,
            I => \N__26857\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26862\,
            I => \N__26854\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26849\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26849\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26846\
        );

    \I__4163\ : Span4Mux_h
    port map (
            O => \N__26854\,
            I => \N__26843\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26840\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26846\,
            I => \N__26837\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__26843\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__4159\ : Odrv12
    port map (
            O => \N__26840\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__26837\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26827\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26827\,
            I => \N__26824\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__26821\,
            I => \N__26817\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26814\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__26817\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26814\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__26809\,
            I => \N__26806\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26800\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26800\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26800\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26794\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26783\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26783\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26780\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__26788\,
            I => \N__26777\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26774\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26780\,
            I => \N__26771\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__26777\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__26774\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__26771\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26761\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__4133\ : Span4Mux_v
    port map (
            O => \N__26758\,
            I => \N__26755\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__26755\,
            I => \N__26751\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26748\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__26751\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26748\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26737\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26737\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__26737\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26731\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26728\
        );

    \I__4123\ : Span4Mux_h
    port map (
            O => \N__26728\,
            I => \N__26723\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26720\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26717\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__26723\,
            I => \N__26714\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__26720\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26717\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__26714\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26702\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26699\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26696\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26693\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26690\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26696\,
            I => \N__26687\
        );

    \I__4110\ : Span4Mux_h
    port map (
            O => \N__26693\,
            I => \N__26683\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__26690\,
            I => \N__26678\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__26687\,
            I => \N__26678\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26675\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__26683\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__26678\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26675\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26659\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26659\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26659\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26656\,
            I => \N__26653\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26653\,
            I => \N__26649\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26646\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__26649\,
            I => \N__26640\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26646\,
            I => \N__26640\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26637\
        );

    \I__4093\ : Span4Mux_h
    port map (
            O => \N__26640\,
            I => \N__26634\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26637\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__26634\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26629\,
            I => \N__26625\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26622\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26617\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26622\,
            I => \N__26617\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__26617\,
            I => \N__26612\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26607\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26607\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__26612\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26607\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26598\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26595\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__26598\,
            I => \N__26590\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26587\
        );

    \I__4077\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26584\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26581\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__26590\,
            I => \N__26578\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__26587\,
            I => \N__26575\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26570\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26570\
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__26578\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__26575\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__26570\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26560\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26560\,
            I => \N__26556\
        );

    \I__4066\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26552\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__26556\,
            I => \N__26549\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26546\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26552\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__26549\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__26546\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4060\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26534\
        );

    \I__4059\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26531\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26528\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26534\,
            I => \N__26525\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__26531\,
            I => \N__26520\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__26528\,
            I => \N__26520\
        );

    \I__4054\ : Span4Mux_v
    port map (
            O => \N__26525\,
            I => \N__26514\
        );

    \I__4053\ : Span4Mux_v
    port map (
            O => \N__26520\,
            I => \N__26514\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26511\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__26514\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__26511\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4049\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26499\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26496\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__26499\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26496\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26486\
        );

    \I__4043\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26481\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26481\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26475\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26481\,
            I => \N__26475\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__26480\,
            I => \N__26472\
        );

    \I__4038\ : Span4Mux_v
    port map (
            O => \N__26475\,
            I => \N__26469\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26466\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__26469\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__26466\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26456\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26453\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26449\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26456\,
            I => \N__26446\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__26453\,
            I => \N__26443\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26440\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26437\
        );

    \I__4027\ : Span12Mux_h
    port map (
            O => \N__26446\,
            I => \N__26434\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__26443\,
            I => \N__26431\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26428\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__26437\,
            I => \N__26425\
        );

    \I__4023\ : Odrv12
    port map (
            O => \N__26434\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__26431\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__26428\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__26425\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26413\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__26410\,
            I => \N__26406\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26402\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__26406\,
            I => \N__26399\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26396\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__26402\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__26399\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__26396\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__26389\,
            I => \N__26384\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26381\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26375\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26375\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26381\,
            I => \N__26372\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26369\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26366\
        );

    \I__4003\ : Span4Mux_h
    port map (
            O => \N__26372\,
            I => \N__26363\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__26369\,
            I => \N__26360\
        );

    \I__4001\ : Span4Mux_h
    port map (
            O => \N__26366\,
            I => \N__26357\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__26363\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__26360\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__26357\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3997\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26346\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26343\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26337\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26337\
        );

    \I__3993\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26334\
        );

    \I__3992\ : Span12Mux_s11_v
    port map (
            O => \N__26337\,
            I => \N__26331\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__26334\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__3990\ : Odrv12
    port map (
            O => \N__26331\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26323\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26317\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26312\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26312\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26309\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__26317\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26312\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__26309\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__3981\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26299\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26295\
        );

    \I__3979\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26292\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__26295\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__26292\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26281\
        );

    \I__3975\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26276\
        );

    \I__3974\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26276\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26273\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26281\,
            I => \N__26268\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26268\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__26273\,
            I => \N__26265\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__26268\,
            I => \N__26260\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__26265\,
            I => \N__26260\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__26260\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26253\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26250\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__26253\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26250\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \N__26242\
        );

    \I__3961\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26239\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26236\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26236\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26226\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26226\
        );

    \I__3956\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26223\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__26226\,
            I => \N__26220\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__26223\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__26220\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \N__26212\
        );

    \I__3951\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26205\
        );

    \I__3950\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26205\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26202\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26205\,
            I => \N__26199\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__26202\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__3946\ : Odrv12
    port map (
            O => \N__26199\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26191\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__26188\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__26182\,
            I => \N__26179\
        );

    \I__3940\ : Span4Mux_h
    port map (
            O => \N__26179\,
            I => \N__26176\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__26176\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26170\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__26170\,
            I => \N__26166\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26163\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26159\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26156\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26153\
        );

    \I__3932\ : Span4Mux_h
    port map (
            O => \N__26159\,
            I => \N__26148\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__26156\,
            I => \N__26148\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__26153\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__26148\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26138\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26135\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26132\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26128\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26125\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26122\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__26131\,
            I => \N__26119\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__26128\,
            I => \N__26114\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__26125\,
            I => \N__26114\
        );

    \I__3919\ : Span4Mux_h
    port map (
            O => \N__26122\,
            I => \N__26111\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26108\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__26114\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__26111\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__26108\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__26101\,
            I => \N__26098\
        );

    \I__3913\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26092\
        );

    \I__3912\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26092\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__26092\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__26089\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26080\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26080\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__26080\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__3906\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26073\
        );

    \I__3905\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26069\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26073\,
            I => \N__26065\
        );

    \I__3903\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26062\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__26069\,
            I => \N__26059\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26056\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__26065\,
            I => \N__26053\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26050\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__26059\,
            I => \N__26045\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__26056\,
            I => \N__26045\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__26053\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3895\ : Odrv12
    port map (
            O => \N__26050\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__26045\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3893\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__26035\,
            I => \N__26031\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26034\,
            I => \N__26027\
        );

    \I__3890\ : Span4Mux_v
    port map (
            O => \N__26031\,
            I => \N__26024\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26021\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__26027\,
            I => \N__26018\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__26024\,
            I => \N__26015\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26021\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__26018\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__26015\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3883\ : InMux
    port map (
            O => \N__26008\,
            I => \N__26005\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__26005\,
            I => \N__26002\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__26002\,
            I => \N__25998\
        );

    \I__3880\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25995\
        );

    \I__3879\ : Span4Mux_v
    port map (
            O => \N__25998\,
            I => \N__25989\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25995\,
            I => \N__25989\
        );

    \I__3877\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25986\
        );

    \I__3876\ : Span4Mux_h
    port map (
            O => \N__25989\,
            I => \N__25983\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25986\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__25983\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__25978\,
            I => \N__25975\
        );

    \I__3872\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__25972\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3870\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25966\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__25966\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__25963\,
            I => \N__25960\
        );

    \I__3867\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25957\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__25957\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25947\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25947\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25944\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25941\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25944\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25941\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__25936\,
            I => \N__25933\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25926\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25926\
        );

    \I__3856\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25923\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25926\,
            I => \N__25920\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25923\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__25920\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__3852\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25912\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__25912\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__25909\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25903\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25897\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25897\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__25897\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__25894\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25885\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25885\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25885\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__25882\,
            I => \N__25879\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25876\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25876\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25869\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25866\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25869\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25866\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25857\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25854\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25857\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25854\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__25849\,
            I => \N__25845\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__25848\,
            I => \N__25842\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25839\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25835\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__25839\,
            I => \N__25832\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25829\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__25835\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__25832\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__25829\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__25822\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__3818\ : Span12Mux_s11_h
    port map (
            O => \N__25813\,
            I => \N__25810\
        );

    \I__3817\ : Odrv12
    port map (
            O => \N__25810\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__3816\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25804\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25804\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__25801\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__25798\,
            I => \N__25795\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25792\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__25792\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25786\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25780\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__25780\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25774\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__3804\ : Odrv12
    port map (
            O => \N__25771\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__3801\ : Odrv12
    port map (
            O => \N__25762\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25755\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25752\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25755\,
            I => \N__25749\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25746\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__25749\,
            I => \N__25739\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__25746\,
            I => \N__25739\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25734\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25734\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__25739\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25734\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25723\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__3787\ : Span12Mux_h
    port map (
            O => \N__25720\,
            I => \N__25717\
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__25717\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__25714\,
            I => \N__25711\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25708\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__25705\,
            I => \N__25702\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__25699\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25690\,
            I => \N__25687\
        );

    \I__3776\ : Sp12to4
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__3775\ : Odrv12
    port map (
            O => \N__25684\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__25681\,
            I => \N__25678\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25675\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__25666\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25654\
        );

    \I__3765\ : Span4Mux_v
    port map (
            O => \N__25654\,
            I => \N__25651\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__25648\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \N__25642\
        );

    \I__3761\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__25636\,
            I => \N__25633\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__25633\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25624\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25624\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25624\,
            I => \N__25619\
        );

    \I__3754\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25614\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25614\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__25619\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25614\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25606\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__25606\,
            I => \N__25603\
        );

    \I__3748\ : Odrv12
    port map (
            O => \N__25603\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25597\,
            I => \N__25594\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__25591\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25585\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__25582\,
            I => \N__25579\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__25579\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__25576\,
            I => \N__25573\
        );

    \I__3738\ : InMux
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__25570\,
            I => \N__25567\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__25567\,
            I => \N__25564\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__25564\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25558\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25558\,
            I => \N__25555\
        );

    \I__3732\ : Span4Mux_v
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__25552\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25546\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25546\,
            I => \N__25543\
        );

    \I__3728\ : Span4Mux_v
    port map (
            O => \N__25543\,
            I => \N__25540\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__25540\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__3726\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25534\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__25534\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__25531\,
            I => \N__25528\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25525\,
            I => \N__25522\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__25522\,
            I => \N__25519\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__25519\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25513\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25513\,
            I => \N__25510\
        );

    \I__3717\ : Odrv4
    port map (
            O => \N__25510\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25504\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25501\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__25501\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25495\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25492\
        );

    \I__3711\ : Span4Mux_v
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__25489\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__25486\,
            I => \N__25483\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25480\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25477\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__25477\,
            I => \N__25474\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__25474\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \N__25468\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25465\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25465\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__25462\,
            I => \N__25459\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25456\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__25456\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__25453\,
            I => \N__25450\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__25447\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__25444\,
            I => \N__25441\
        );

    \I__3694\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__25438\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__25432\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__25429\,
            I => \N__25426\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__3687\ : Span4Mux_v
    port map (
            O => \N__25420\,
            I => \N__25417\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__25417\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25411\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__25411\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__25402\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__3680\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__3678\ : Odrv12
    port map (
            O => \N__25393\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25387\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__25387\,
            I => \N__25384\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__25384\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__3674\ : InMux
    port map (
            O => \N__25381\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__25378\,
            I => \N__25353\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25342\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25342\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25327\
        );

    \I__3669\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25327\
        );

    \I__3668\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25327\
        );

    \I__3667\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25327\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25327\
        );

    \I__3665\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25327\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25327\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25310\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25310\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25310\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25310\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25310\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25310\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25310\
        );

    \I__3656\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25310\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25299\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25299\
        );

    \I__3653\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25299\
        );

    \I__3652\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25299\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25299\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25296\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25280\
        );

    \I__3648\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25280\
        );

    \I__3647\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25280\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25280\
        );

    \I__3645\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25280\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25280\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25271\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25327\,
            I => \N__25271\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__25310\,
            I => \N__25271\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25299\,
            I => \N__25271\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__25296\,
            I => \N__25268\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25263\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25263\
        );

    \I__3636\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25260\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25255\
        );

    \I__3634\ : Span4Mux_v
    port map (
            O => \N__25271\,
            I => \N__25255\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__25268\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__25263\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25260\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__25255\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25246\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25243\,
            I => \N__25240\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__25240\,
            I => \N__25237\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__25237\,
            I => \N__25234\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__25234\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__25228\,
            I => \N__25225\
        );

    \I__3622\ : Odrv4
    port map (
            O => \N__25225\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25219\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__25219\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__3618\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25210\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__25210\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__25207\,
            I => \N__25204\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25201\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__25201\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__25198\,
            I => \N__25195\
        );

    \I__3612\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25192\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__25192\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__25183\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25177\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25174\
        );

    \I__3605\ : Span4Mux_h
    port map (
            O => \N__25174\,
            I => \N__25171\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__25171\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25168\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25162\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__25162\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25159\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25153\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25150\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__25150\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25147\,
            I => \bfn_10_17_0_\
        );

    \I__3595\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__3593\ : Odrv12
    port map (
            O => \N__25138\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25135\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__25126\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25123\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25117\,
            I => \N__25114\
        );

    \I__3585\ : Odrv12
    port map (
            O => \N__25114\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25111\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25105\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__25102\,
            I => \N__25099\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__25099\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__3579\ : InMux
    port map (
            O => \N__25096\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__3578\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25090\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__25090\,
            I => \N__25087\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__25087\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__3575\ : InMux
    port map (
            O => \N__25084\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__3574\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25078\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25078\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__3572\ : InMux
    port map (
            O => \N__25075\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__3571\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25069\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__25069\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25066\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__3568\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25060\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25060\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__3566\ : InMux
    port map (
            O => \N__25057\,
            I => \bfn_10_16_0_\
        );

    \I__3565\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25051\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25051\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__3563\ : InMux
    port map (
            O => \N__25048\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25042\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25039\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25033\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__25030\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__3556\ : InMux
    port map (
            O => \N__25027\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25021\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__25018\,
            I => \N__25015\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__25015\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25012\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__25003\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25000\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24994\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__24994\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24991\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24985\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__24985\,
            I => \N__24982\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__24982\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24979\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24973\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__24973\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__3537\ : InMux
    port map (
            O => \N__24970\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__24964\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24961\,
            I => \bfn_10_15_0_\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24955\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__24955\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24952\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24946\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__3528\ : Span4Mux_v
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__24940\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24937\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24931\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__24928\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24925\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24919\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24916\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24916\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24913\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24907\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24907\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__3515\ : InMux
    port map (
            O => \N__24904\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24896\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24893\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24890\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24887\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24893\,
            I => \N__24884\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24890\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__3508\ : Odrv12
    port map (
            O => \N__24887\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__24884\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24872\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24869\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24866\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24863\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24869\,
            I => \N__24860\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__24866\,
            I => \N__24857\
        );

    \I__3500\ : Span4Mux_v
    port map (
            O => \N__24863\,
            I => \N__24853\
        );

    \I__3499\ : Span4Mux_v
    port map (
            O => \N__24860\,
            I => \N__24848\
        );

    \I__3498\ : Span4Mux_v
    port map (
            O => \N__24857\,
            I => \N__24848\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24845\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__24853\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__24848\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24845\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24833\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24828\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24836\,
            I => \N__24828\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24824\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24828\,
            I => \N__24821\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24818\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__24824\,
            I => \N__24813\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__24821\,
            I => \N__24813\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24818\,
            I => \N__24810\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__24813\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__24810\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24798\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24795\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__24798\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24795\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24787\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24784\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24778\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24778\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24775\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \N__24765\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24760\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24760\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24760\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24748\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24748\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24748\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__3459\ : Span4Mux_h
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__24733\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__24730\,
            I => \N__24726\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24721\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24721\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24718\
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__24718\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__24715\,
            I => \N__24711\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24705\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24705\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24702\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24705\,
            I => \N__24699\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24702\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24699\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24687\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24687\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24684\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24681\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__24684\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__24681\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24673\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__24670\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__24667\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24658\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24658\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__24655\,
            I => \N__24652\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24649\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24646\
        );

    \I__3429\ : Odrv12
    port map (
            O => \N__24646\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24637\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__24634\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__3421\ : Odrv12
    port map (
            O => \N__24622\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24619\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24610\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__24610\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__24607\,
            I => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24595\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__24595\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__24592\,
            I => \N__24587\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24584\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24579\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24579\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24584\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24579\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24569\
        );

    \I__3404\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24564\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24564\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__24569\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__24564\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24556\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24556\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24550\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__24541\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24534\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24531\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__24534\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24531\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__24526\,
            I => \N__24523\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24520\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__24517\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24511\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__24511\,
            I => \N__24508\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__24505\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__3381\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24498\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24495\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__24498\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24495\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__24490\,
            I => \N__24487\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24484\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__24475\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24468\
        );

    \I__3370\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24465\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__24468\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__24465\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__24460\,
            I => \N__24457\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24454\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__24454\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__24448\,
            I => \N__24445\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__24445\,
            I => \N__24442\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__24442\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24439\,
            I => \N__24436\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24433\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24433\,
            I => \N__24430\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__24427\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__3355\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24418\
        );

    \I__3353\ : Span4Mux_h
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__24415\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__3350\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24406\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24406\,
            I => \N__24403\
        );

    \I__3348\ : Span4Mux_h
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__24400\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24394\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__24391\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24382\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__3340\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24373\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__24373\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3337\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24366\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24363\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__24366\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__24363\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24352\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24345\
        );

    \I__3329\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24342\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24345\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__24342\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24334\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24334\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24327\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24324\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24327\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24324\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__24319\,
            I => \N__24316\
        );

    \I__3319\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24313\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__24313\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3317\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24306\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24303\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__24306\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__24303\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24295\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__24295\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24288\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24285\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__24288\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24277\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__24277\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24270\
        );

    \I__3304\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24267\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__24270\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__24267\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24252\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24249\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24252\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24249\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__24244\,
            I => \N__24241\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24238\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__24238\,
            I => \N__24235\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__24235\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24228\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24225\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24228\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24225\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__24220\,
            I => \N__24217\
        );

    \I__3286\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24214\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24211\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__24211\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__24208\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__3281\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24199\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24199\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__24196\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24190\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24190\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24178\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24175\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__24175\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__3271\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24168\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24165\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__24168\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__24165\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__24160\,
            I => \N__24157\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24154\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__24154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24147\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24144\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__24147\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__24144\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24136\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__24136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3258\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24130\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24127\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__24127\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24120\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24117\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__24120\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24117\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__24112\,
            I => \N__24109\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24106\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__24106\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24099\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24096\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__24099\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24096\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__24091\,
            I => \N__24087\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24083\
        );

    \I__3242\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24080\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24077\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24083\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__24080\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__24077\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24070\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24067\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__3235\ : IoInMux
    port map (
            O => \N__24064\,
            I => \N__24061\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__3233\ : Span4Mux_s1_v
    port map (
            O => \N__24058\,
            I => \N__24055\
        );

    \I__3232\ : Span4Mux_v
    port map (
            O => \N__24055\,
            I => \N__24051\
        );

    \I__3231\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24048\
        );

    \I__3230\ : Sp12to4
    port map (
            O => \N__24051\,
            I => \N__24044\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24041\
        );

    \I__3228\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24038\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__24044\,
            I => s1_phy_c
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__24041\,
            I => s1_phy_c
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__24038\,
            I => s1_phy_c
        );

    \I__3224\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24026\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24021\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24021\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__24026\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__24021\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3219\ : InMux
    port map (
            O => \N__24016\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__24013\,
            I => \N__24009\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24005\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24009\,
            I => \N__24002\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23999\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__24005\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__24002\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23999\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23992\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__23989\,
            I => \N__23984\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__23988\,
            I => \N__23981\
        );

    \I__3208\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23978\
        );

    \I__3207\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23973\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23973\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__23978\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__23973\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23968\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23960\
        );

    \I__3201\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23955\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23955\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23960\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23955\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23950\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__3196\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23942\
        );

    \I__3195\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23937\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23937\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23942\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23937\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23932\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__23929\,
            I => \N__23925\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__23928\,
            I => \N__23921\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23918\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23915\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23912\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23918\,
            I => \N__23909\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__23915\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__23912\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__23909\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__3181\ : InMux
    port map (
            O => \N__23902\,
            I => \bfn_9_23_0_\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__23899\,
            I => \N__23895\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__23898\,
            I => \N__23891\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23895\,
            I => \N__23888\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23885\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23882\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23879\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23885\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__23882\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__23879\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23872\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23865\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23862\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23865\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23862\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__23857\,
            I => \N__23853\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23849\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23846\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23843\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23849\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23846\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__23843\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23836\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__23833\,
            I => \N__23829\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23825\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23822\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23819\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23825\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__23822\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23819\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23812\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23804\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23799\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23799\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23804\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23799\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23794\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__23791\,
            I => \N__23787\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23783\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23780\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23777\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__23783\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23780\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23777\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23770\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__23767\,
            I => \N__23762\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__23766\,
            I => \N__23759\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23756\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23751\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23751\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23756\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23751\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23746\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23733\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23733\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23738\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23733\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23728\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23720\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23724\,
            I => \N__23715\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23715\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23720\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23715\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23710\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__23707\,
            I => \N__23703\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__23706\,
            I => \N__23699\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23696\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23693\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23690\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23687\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23693\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__23690\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__23687\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23680\,
            I => \bfn_9_22_0_\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23673\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23670\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23666\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23663\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23660\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__23666\,
            I => \N__23657\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23654\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23660\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__23657\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__23654\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23647\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__23644\,
            I => \N__23640\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23636\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23633\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23630\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23636\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23633\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__23630\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3088\ : InMux
    port map (
            O => \N__23623\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__23620\,
            I => \N__23615\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__23619\,
            I => \N__23612\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23604\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23604\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23609\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__23604\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23599\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__23596\,
            I => \N__23592\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23583\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23583\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23580\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23577\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23580\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__23577\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23572\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__23569\,
            I => \N__23565\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23561\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23558\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23555\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__23558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__23555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23548\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23541\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23537\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23534\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23531\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__23537\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__23534\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23531\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23524\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23516\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23511\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23511\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23516\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__23511\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3049\ : InMux
    port map (
            O => \N__23506\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23498\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23493\
        );

    \I__3046\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23493\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23498\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__23493\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3043\ : InMux
    port map (
            O => \N__23488\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23482\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23478\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__23481\,
            I => \N__23474\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23471\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23468\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23465\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__23471\,
            I => \N__23462\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__23468\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__23465\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__23462\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3032\ : InMux
    port map (
            O => \N__23455\,
            I => \bfn_9_21_0_\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__23452\,
            I => \N__23448\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__23451\,
            I => \N__23444\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23441\
        );

    \I__3028\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23438\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23435\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23432\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__23438\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23435\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__23432\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23425\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23422\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23419\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23413\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__23413\,
            I => \N__23410\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__23410\,
            I => \N__23407\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__23407\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23401\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23401\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__23398\,
            I => \N__23395\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__23392\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23386\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__23383\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23377\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__23377\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__23371\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23365\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__23365\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23359\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23359\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__2999\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23353\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23353\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__2997\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23347\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23347\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23341\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23341\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__2993\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23335\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__23335\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23329\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23329\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23323\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__23323\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__2987\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23317\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__23317\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23311\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23308\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__23305\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__2981\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23296\
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__23296\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__23293\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__23290\,
            I => \N__23285\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23282\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23279\
        );

    \I__2974\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23276\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23282\,
            I => \current_shift_inst.N_1306_i\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__23279\,
            I => \current_shift_inst.N_1306_i\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__23276\,
            I => \current_shift_inst.N_1306_i\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23266\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__23266\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23260\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__23260\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23254\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__23254\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23248\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23248\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__23245\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23241\,
            I => \N__23236\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__23236\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23228\
        );

    \I__2957\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23223\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23223\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23228\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__23223\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__23218\,
            I => \N__23214\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__23217\,
            I => \N__23211\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23206\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23206\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__23200\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23190\
        );

    \I__2945\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23190\
        );

    \I__2944\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23187\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23190\,
            I => \N__23184\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23187\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__23184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__23179\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23170\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__23167\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \N__23161\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__23158\,
            I => \N__23155\
        );

    \I__2932\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__23152\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23146\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23146\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23140\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23137\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23134\,
            I => \bfn_9_10_0_\
        );

    \I__2924\ : InMux
    port map (
            O => \N__23131\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__2923\ : InMux
    port map (
            O => \N__23128\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23125\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__2921\ : InMux
    port map (
            O => \N__23122\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__23119\,
            I => \N__23115\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23112\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23109\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__23112\,
            I => \N__23103\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23103\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23100\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__23103\,
            I => \N__23097\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__23100\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__23097\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__2911\ : InMux
    port map (
            O => \N__23092\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23089\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \N__23082\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23076\
        );

    \I__2907\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23076\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23073\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23076\,
            I => \N__23070\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23073\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__2903\ : Odrv12
    port map (
            O => \N__23070\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23065\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__23062\,
            I => \N__23057\
        );

    \I__2900\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23054\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23051\
        );

    \I__2898\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23048\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23045\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__23051\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23048\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__23045\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23038\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23029\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__23029\,
            I => \N__23024\
        );

    \I__2889\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23021\
        );

    \I__2888\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23018\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__23024\,
            I => \N__23015\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__23012\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__23018\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__23015\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__23012\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23005\,
            I => \bfn_9_9_0_\
        );

    \I__2881\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22997\
        );

    \I__2880\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22992\
        );

    \I__2879\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22992\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__22997\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__22992\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22987\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22979\
        );

    \I__2874\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22974\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22974\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__22979\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22974\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22969\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22966\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22963\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22960\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22957\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__2865\ : InMux
    port map (
            O => \N__22954\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22951\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22948\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22945\,
            I => \bfn_9_8_0_\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22942\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22939\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22936\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22933\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22930\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22927\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22900\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22900\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22900\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22900\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22891\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22891\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22891\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22891\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22868\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22868\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22868\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22868\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22859\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22859\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22859\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22859\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22854\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22891\,
            I => \N__22854\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22849\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22849\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22840\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22840\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22840\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22840\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22884\,
            I => \N__22831\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22831\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22831\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22831\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22822\
        );

    \I__2826\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22822\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22822\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22877\,
            I => \N__22822\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22817\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22817\
        );

    \I__2821\ : Span4Mux_h
    port map (
            O => \N__22854\,
            I => \N__22814\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__22849\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22840\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22831\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22822\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__22817\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__22814\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22801\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__2813\ : CEMux
    port map (
            O => \N__22798\,
            I => \N__22794\
        );

    \I__2812\ : CEMux
    port map (
            O => \N__22797\,
            I => \N__22791\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22788\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22785\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__22788\,
            I => \N__22780\
        );

    \I__2808\ : Span12Mux_h
    port map (
            O => \N__22785\,
            I => \N__22777\
        );

    \I__2807\ : CEMux
    port map (
            O => \N__22784\,
            I => \N__22774\
        );

    \I__2806\ : CEMux
    port map (
            O => \N__22783\,
            I => \N__22771\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__22780\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__22777\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22774\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22771\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__22762\,
            I => \N__22757\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22753\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22748\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22748\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22745\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22753\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22748\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22745\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22738\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__2792\ : InMux
    port map (
            O => \N__22735\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__2791\ : InMux
    port map (
            O => \N__22732\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22729\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22726\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22723\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22720\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22717\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__2785\ : InMux
    port map (
            O => \N__22714\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22711\,
            I => \bfn_8_24_0_\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22708\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__2782\ : InMux
    port map (
            O => \N__22705\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22702\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__2780\ : InMux
    port map (
            O => \N__22699\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22696\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22693\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22690\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22687\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22684\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22681\,
            I => \bfn_8_23_0_\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22678\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22675\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22672\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22669\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__2769\ : InMux
    port map (
            O => \N__22666\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22663\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22660\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22657\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22654\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__2764\ : InMux
    port map (
            O => \N__22651\,
            I => \bfn_8_22_0_\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22648\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__2762\ : CEMux
    port map (
            O => \N__22645\,
            I => \N__22639\
        );

    \I__2761\ : CEMux
    port map (
            O => \N__22644\,
            I => \N__22636\
        );

    \I__2760\ : CEMux
    port map (
            O => \N__22643\,
            I => \N__22633\
        );

    \I__2759\ : CEMux
    port map (
            O => \N__22642\,
            I => \N__22630\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22624\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__22636\,
            I => \N__22624\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22633\,
            I => \N__22621\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22630\,
            I => \N__22618\
        );

    \I__2754\ : CEMux
    port map (
            O => \N__22629\,
            I => \N__22615\
        );

    \I__2753\ : Span4Mux_v
    port map (
            O => \N__22624\,
            I => \N__22606\
        );

    \I__2752\ : Span4Mux_v
    port map (
            O => \N__22621\,
            I => \N__22606\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__22618\,
            I => \N__22606\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22606\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__22606\,
            I => \N__22603\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__22600\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__22597\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22591\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__22591\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__22588\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22585\,
            I => \bfn_8_21_0_\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22579\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22552\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22552\
        );

    \I__2737\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22552\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22552\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22533\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22533\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22533\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22533\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22520\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22520\
        );

    \I__2729\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22520\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22520\
        );

    \I__2727\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22511\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22511\
        );

    \I__2725\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22511\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22511\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__22552\,
            I => \N__22508\
        );

    \I__2722\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22499\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22499\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22499\
        );

    \I__2719\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22499\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22494\
        );

    \I__2717\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22494\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22485\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22485\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22485\
        );

    \I__2713\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22485\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22482\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22473\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22473\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22473\
        );

    \I__2708\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22473\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22470\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22463\
        );

    \I__2705\ : Span4Mux_h
    port map (
            O => \N__22508\,
            I => \N__22463\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22463\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22454\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__22485\,
            I => \N__22454\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__22482\,
            I => \N__22454\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22473\,
            I => \N__22454\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__22470\,
            I => \N__22449\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__22463\,
            I => \N__22449\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__22454\,
            I => \N__22446\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__22449\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__22446\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__22435\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__2691\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__22426\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__22417\,
            I => \N__22414\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__22414\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__2684\ : CEMux
    port map (
            O => \N__22411\,
            I => \N__22406\
        );

    \I__2683\ : CEMux
    port map (
            O => \N__22410\,
            I => \N__22403\
        );

    \I__2682\ : CEMux
    port map (
            O => \N__22409\,
            I => \N__22400\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22396\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22403\,
            I => \N__22393\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22390\
        );

    \I__2678\ : CEMux
    port map (
            O => \N__22399\,
            I => \N__22387\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__22396\,
            I => \N__22384\
        );

    \I__2676\ : Span4Mux_v
    port map (
            O => \N__22393\,
            I => \N__22379\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__22390\,
            I => \N__22379\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22376\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__22384\,
            I => \N__22371\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__22379\,
            I => \N__22371\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__22376\,
            I => \N__22368\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__22371\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__22368\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__2668\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22357\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22357\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22352\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22347\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22347\
        );

    \I__2663\ : Span12Mux_v
    port map (
            O => \N__22352\,
            I => \N__22344\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__22347\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__22344\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22326\
        );

    \I__2658\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22326\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22326\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22323\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__22326\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22323\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22309\
        );

    \I__2652\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22309\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22309\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__22309\,
            I => \N__22306\
        );

    \I__2649\ : Span12Mux_v
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__2648\ : Odrv12
    port map (
            O => \N__22303\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__2647\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22297\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22297\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22294\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__2644\ : InMux
    port map (
            O => \N__22291\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__22285\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__22279\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22270\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__22270\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22263\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22260\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22263\,
            I => \current_shift_inst.control_input_31\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22260\,
            I => \current_shift_inst.control_input_31\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__22252\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__22243\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__22234\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__22228\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22222\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__2620\ : InMux
    port map (
            O => \N__22219\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__2619\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22213\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__22213\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22210\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22204\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22201\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__2613\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22195\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__22195\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22192\,
            I => \bfn_8_16_0_\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22186\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__2608\ : InMux
    port map (
            O => \N__22183\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22177\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22177\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22174\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22168\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__2602\ : InMux
    port map (
            O => \N__22165\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__22159\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22156\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22153\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__22147\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22144\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__2594\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22138\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__22138\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22135\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__22129\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22126\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__22120\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__2586\ : InMux
    port map (
            O => \N__22117\,
            I => \bfn_8_15_0_\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__22111\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22108\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__2582\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__22102\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22099\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__22093\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22090\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22084\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22084\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22081\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22075\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__22075\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22072\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__22066\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__2568\ : InMux
    port map (
            O => \N__22063\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__2567\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__22057\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22054\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__22048\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22045\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__22039\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__2559\ : InMux
    port map (
            O => \N__22036\,
            I => \bfn_8_14_0_\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22030\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__22030\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__2556\ : InMux
    port map (
            O => \N__22027\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__22021\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__2553\ : InMux
    port map (
            O => \N__22018\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22012\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22012\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__2550\ : InMux
    port map (
            O => \N__22009\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__2549\ : InMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22003\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21992\
        );

    \I__2545\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21989\
        );

    \I__2544\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21986\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21983\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__21989\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__21986\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__21983\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21976\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__2538\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21969\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21966\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__21969\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__21966\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__21961\,
            I => \N__21958\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21953\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21950\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21947\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21953\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21950\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21947\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21940\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21933\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21930\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21933\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__21930\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__21925\,
            I => \N__21920\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__21924\,
            I => \N__21917\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21914\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21909\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21909\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__21914\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21909\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21904\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21901\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__21895\,
            I => \current_shift_inst.control_input_1\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21889\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21886\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__21880\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21877\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21871\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21868\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__21865\,
            I => \N__21861\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__21864\,
            I => \N__21858\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21854\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21851\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21848\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21845\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__21851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21848\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__21845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21838\,
            I => \bfn_8_11_0_\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__21835\,
            I => \N__21831\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__21834\,
            I => \N__21828\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21824\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21821\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21818\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21815\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21821\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21818\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21808\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__21805\,
            I => \N__21802\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21797\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21794\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21791\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21797\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21794\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__21791\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21784\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21776\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21771\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21771\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21776\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21771\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21766\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21763\,
            I => \N__21760\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21755\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21752\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21749\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21755\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21752\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21749\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21742\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__21739\,
            I => \N__21734\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__21738\,
            I => \N__21731\
        );

    \I__2458\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21728\
        );

    \I__2457\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21723\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21723\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__21728\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21723\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21718\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21710\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21705\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21705\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21710\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21705\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21700\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21692\
        );

    \I__2445\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21687\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21687\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21692\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21687\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21682\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__21679\,
            I => \N__21675\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__21678\,
            I => \N__21672\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21668\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21665\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21662\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N__21659\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21662\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__21659\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21652\,
            I => \bfn_8_12_0_\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__21649\,
            I => \N__21645\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__21648\,
            I => \N__21642\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21638\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21635\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21632\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21629\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__21635\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__21632\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__21629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21622\,
            I => \bfn_8_10_0_\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21612\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__21615\,
            I => \N__21609\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21605\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21602\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21599\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__21605\,
            I => \N__21596\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21602\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21599\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__21596\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21589\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21578\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21575\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21572\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__21578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__21575\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21572\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21560\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__21564\,
            I => \N__21556\
        );

    \I__2400\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21553\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21550\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21545\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21545\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21553\,
            I => \N__21542\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__21550\,
            I => \N__21539\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__21545\,
            I => \N__21536\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__21542\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__21539\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__21536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21529\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21521\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21516\
        );

    \I__2387\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21516\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21521\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__21516\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21511\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__2382\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21500\
        );

    \I__2381\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21497\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21494\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__21500\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__21497\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21494\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21487\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__21484\,
            I => \N__21479\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__21483\,
            I => \N__21476\
        );

    \I__2373\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21473\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21468\
        );

    \I__2371\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21468\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__21473\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__21468\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21463\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21455\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21450\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21450\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__21455\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__21450\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21445\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21437\
        );

    \I__2360\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21432\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21432\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__21432\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21427\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__21424\,
            I => \N__21420\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21416\
        );

    \I__2353\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21413\
        );

    \I__2352\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21410\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__21416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__21413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__21410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__2347\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21396\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21392\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__21396\,
            I => \N__21389\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21386\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__21392\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__21389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21386\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2340\ : InMux
    port map (
            O => \N__21379\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__2339\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21371\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21366\
        );

    \I__2337\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21366\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__21371\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__21366\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__2334\ : InMux
    port map (
            O => \N__21361\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__21358\,
            I => \N__21355\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21350\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21347\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21344\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__21350\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__21347\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__21344\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__2326\ : InMux
    port map (
            O => \N__21337\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__21334\,
            I => \N__21329\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__21333\,
            I => \N__21326\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21323\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21318\
        );

    \I__2321\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21318\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__21323\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21318\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21313\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__21310\,
            I => \N__21307\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21302\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21299\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21296\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21302\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21299\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21296\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21289\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21281\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21276\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21276\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21281\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21276\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21271\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21263\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21258\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21258\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21263\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__21258\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21253\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21246\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21243\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21246\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__21243\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__21238\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21231\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21228\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21231\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21228\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__21223\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21214\
        );

    \I__2286\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21214\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__21214\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__21211\,
            I => \N__21207\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__21210\,
            I => \N__21204\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21199\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21199\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21196\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__21196\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__2278\ : InMux
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__21190\,
            I => \N__21187\
        );

    \I__2276\ : Span4Mux_s3_h
    port map (
            O => \N__21187\,
            I => \N__21183\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21180\
        );

    \I__2274\ : Span4Mux_h
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__21180\,
            I => \N__21174\
        );

    \I__2272\ : Sp12to4
    port map (
            O => \N__21177\,
            I => \N__21171\
        );

    \I__2271\ : Odrv12
    port map (
            O => \N__21174\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__21171\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21158\
        );

    \I__2268\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21158\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21155\
        );

    \I__2266\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21152\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21158\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__21155\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21152\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__2262\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__2261\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21134\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21134\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21131\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21139\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__21134\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21131\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__2255\ : IoInMux
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21118\
        );

    \I__2253\ : Span4Mux_s0_v
    port map (
            O => \N__21118\,
            I => \N__21115\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__21115\,
            I => \N__21112\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__21112\,
            I => \N__21109\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__21109\,
            I => \current_shift_inst.timer_s1.N_161_i\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__21106\,
            I => \N__21103\
        );

    \I__2248\ : GlobalMux
    port map (
            O => \N__21103\,
            I => \N__21100\
        );

    \I__2247\ : gio2CtrlBuf
    port map (
            O => \N__21100\,
            I => delay_hc_input_c_g
        );

    \I__2246\ : InMux
    port map (
            O => \N__21097\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21094\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21091\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__2243\ : InMux
    port map (
            O => \N__21088\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21085\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__2241\ : InMux
    port map (
            O => \N__21082\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21076\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21073\
        );

    \I__2238\ : Span4Mux_s3_h
    port map (
            O => \N__21073\,
            I => \N__21070\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__21070\,
            I => \N__21067\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__21067\,
            I => \N__21063\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21060\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__21063\,
            I => \N__21057\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21060\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__21057\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21052\,
            I => \N__21049\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21049\,
            I => \N__21045\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21042\
        );

    \I__2228\ : Span12Mux_v
    port map (
            O => \N__21045\,
            I => \N__21039\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21042\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__2226\ : Odrv12
    port map (
            O => \N__21039\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21031\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__21031\,
            I => \N__21027\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21024\
        );

    \I__2222\ : Span4Mux_h
    port map (
            O => \N__21027\,
            I => \N__21021\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__21024\,
            I => \N__21018\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__21021\,
            I => \N__21015\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__21018\,
            I => \N__21010\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__21015\,
            I => \N__21010\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__21010\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__2216\ : InMux
    port map (
            O => \N__21007\,
            I => \N__21003\
        );

    \I__2215\ : InMux
    port map (
            O => \N__21006\,
            I => \N__21000\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20997\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__21000\,
            I => \N__20994\
        );

    \I__2212\ : Span12Mux_s7_h
    port map (
            O => \N__20997\,
            I => \N__20991\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__20994\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__20991\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20986\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20983\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20980\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20977\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__2205\ : InMux
    port map (
            O => \N__20974\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20971\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20968\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20965\,
            I => \bfn_7_17_0_\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20962\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20959\,
            I => \bfn_7_15_0_\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20956\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20953\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20950\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20947\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20944\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20941\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20938\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20935\,
            I => \bfn_7_16_0_\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20932\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20926\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__20926\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20923\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20920\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20917\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20914\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20911\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20908\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20905\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20902\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__2180\ : InMux
    port map (
            O => \N__20899\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20896\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20893\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20890\,
            I => \bfn_7_13_0_\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20887\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20884\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20881\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20878\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20875\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20872\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20869\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20866\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20863\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20860\,
            I => \bfn_7_12_0_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20857\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20854\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20851\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20848\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20845\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20842\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20839\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20836\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20833\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20830\,
            I => \bfn_7_11_0_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20827\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20824\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20818\,
            I => \N__20814\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20810\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__20814\,
            I => \N__20807\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20804\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20810\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__20807\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20804\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__20797\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20791\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__20791\,
            I => \N__20788\
        );

    \I__2143\ : Odrv12
    port map (
            O => \N__20788\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20785\,
            I => \bfn_7_10_0_\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20782\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20773\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20773\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20773\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__20770\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20764\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20764\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20758\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20748\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20745\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20748\,
            I => \N__20740\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__20745\,
            I => \N__20740\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__20740\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__20737\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20731\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20725\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20725\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__20722\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__20719\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20713\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__20704\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20698\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__20695\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__20692\,
            I => \N__20682\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__20691\,
            I => \N__20679\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__20690\,
            I => \N__20667\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__20689\,
            I => \N__20664\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__20688\,
            I => \N__20661\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__20687\,
            I => \N__20657\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20638\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20638\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20638\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20638\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20638\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20633\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20633\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20624\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20624\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20624\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20624\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__20671\,
            I => \N__20620\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__20670\,
            I => \N__20617\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20606\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20606\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20606\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20606\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20599\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20599\
        );

    \I__2086\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20599\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20594\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20583\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20583\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20583\
        );

    \I__2081\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20583\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20583\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20580\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20575\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20575\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20572\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20563\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20563\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20563\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20563\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20558\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20558\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20555\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20552\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20594\,
            I => \N__20547\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20583\,
            I => \N__20547\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__20580\,
            I => \N__20542\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__20575\,
            I => \N__20542\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20572\,
            I => \N__20535\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20535\
        );

    \I__2061\ : Sp12to4
    port map (
            O => \N__20558\,
            I => \N__20535\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20528\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20528\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__20547\,
            I => \N__20528\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__20542\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2056\ : Odrv12
    port map (
            O => \N__20535\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__20528\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20518\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__20515\,
            I => \N__20512\
        );

    \I__2051\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20506\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__20506\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20497\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__20497\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__2044\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20488\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20485\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__20482\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20473\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__20467\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20455\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__2028\ : Span4Mux_h
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__20440\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__20437\,
            I => \N__20414\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__20436\,
            I => \N__20411\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__20435\,
            I => \N__20408\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__20434\,
            I => \N__20405\
        );

    \I__2022\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20395\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20386\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20386\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20386\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20386\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__20428\,
            I => \N__20382\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__20427\,
            I => \N__20379\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__20426\,
            I => \N__20374\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__20425\,
            I => \N__20371\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20364\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20364\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20364\
        );

    \I__2010\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20355\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20355\
        );

    \I__2008\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20355\
        );

    \I__2007\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20355\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20352\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20349\
        );

    \I__2004\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20338\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20338\
        );

    \I__2002\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20338\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20338\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20338\
        );

    \I__1999\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20327\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20327\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20400\,
            I => \N__20327\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20327\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20327\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20395\,
            I => \N__20324\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__20386\,
            I => \N__20321\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20318\
        );

    \I__1991\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20313\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20313\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20304\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20304\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20304\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20304\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20364\,
            I => \N__20299\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20299\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20286\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20286\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20338\,
            I => \N__20286\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20286\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__20324\,
            I => \N__20286\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__20321\,
            I => \N__20286\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__20318\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__20313\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20304\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__1974\ : Odrv12
    port map (
            O => \N__20299\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__20286\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20272\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20272\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__20269\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__20263\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__1967\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20257\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__20257\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__20254\,
            I => \N__20251\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20248\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__20248\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__20245\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__20239\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__20236\,
            I => \N__20232\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__20235\,
            I => \N__20229\
        );

    \I__1957\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20226\
        );

    \I__1956\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20223\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20218\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20218\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__20218\,
            I => \N__20215\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__20215\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20209\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__20209\,
            I => \N__20206\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__20206\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__20203\,
            I => \N__20200\
        );

    \I__1947\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__20197\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20191\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20191\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__20185\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__20179\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \N__20173\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20170\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__20170\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__20164\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__20161\,
            I => \N__20158\
        );

    \I__1933\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20155\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__20152\,
            I => \N__20149\
        );

    \I__1930\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__20146\,
            I => \N__20143\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__20143\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20137\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__20137\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1925\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20131\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20131\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20125\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__20125\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__1920\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__20116\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20107\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__20107\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20101\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20101\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__20098\,
            I => \N__20095\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20092\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__20092\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20086\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__20086\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__1907\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20077\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20077\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__1905\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20071\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__20071\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__20068\,
            I => \N__20065\
        );

    \I__1902\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20062\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__20062\,
            I => \N__20059\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__20059\,
            I => \N__20056\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__20056\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1898\ : InMux
    port map (
            O => \N__20053\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__20050\,
            I => \N__20047\
        );

    \I__1896\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20044\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__20044\,
            I => \N__20041\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__20041\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1893\ : InMux
    port map (
            O => \N__20038\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__20035\,
            I => \N__20032\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20029\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__20023\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20020\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__20011\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \N__20005\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19999\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__19996\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19993\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__19990\,
            I => \N__19987\
        );

    \I__1876\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19984\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__19984\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1874\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19978\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__19978\,
            I => \N__19975\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__19975\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__19969\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__1868\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19960\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__19960\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__19951\,
            I => \N_39_i_i\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19942\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__19939\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19936\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__1855\ : Span4Mux_h
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__19921\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19918\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \N__19912\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__19903\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19900\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__1843\ : Span4Mux_h
    port map (
            O => \N__19888\,
            I => \N__19885\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19885\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19882\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__19879\,
            I => \N__19876\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19873\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__19873\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19870\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19861\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19861\,
            I => \N__19858\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__19855\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19852\,
            I => \bfn_2_14_0_\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__19849\,
            I => \N__19846\
        );

    \I__1829\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19843\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__19837\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19834\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__19831\,
            I => \N__19828\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19825\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19822\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__19822\,
            I => \N__19819\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__19819\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19816\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__19813\,
            I => \N__19810\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19807\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19804\
        );

    \I__1815\ : Span4Mux_h
    port map (
            O => \N__19804\,
            I => \N__19801\
        );

    \I__1814\ : Span4Mux_s0_h
    port map (
            O => \N__19801\,
            I => \N__19798\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__19798\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19795\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__19792\,
            I => \N__19789\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19783\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__1807\ : Span4Mux_h
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__19777\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19774\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__1800\ : Span4Mux_h
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__19756\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19753\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__19750\,
            I => \N__19747\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19744\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__19741\,
            I => \N__19738\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__19738\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19735\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__19729\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19726\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1788\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19717\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19717\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19714\,
            I => \bfn_2_13_0_\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19705\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19705\,
            I => \N__19702\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__19702\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19699\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19690\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19687\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19684\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19672\
        );

    \I__1771\ : Span4Mux_h
    port map (
            O => \N__19672\,
            I => \N__19669\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19669\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19666\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19657\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__19654\,
            I => \N__19651\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__19651\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19648\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__19645\,
            I => \N__19642\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19639\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19639\,
            I => \N__19636\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__19633\,
            I => \N__19630\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__19630\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19627\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19618\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19618\,
            I => \N__19615\
        );

    \I__1752\ : Span4Mux_v
    port map (
            O => \N__19615\,
            I => \N__19612\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__19612\,
            I => \N__19609\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__19609\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19606\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__1747\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__19594\,
            I => \N__19591\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__19591\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19588\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19579\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19576\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19573\
        );

    \I__1738\ : Span4Mux_s0_h
    port map (
            O => \N__19573\,
            I => \N__19570\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__19570\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19567\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \N__19561\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19558\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19555\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__19555\,
            I => \N__19552\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__19552\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1730\ : InMux
    port map (
            O => \N__19549\,
            I => \bfn_2_12_0_\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__19546\,
            I => \N__19543\
        );

    \I__1728\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19540\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__19540\,
            I => \N__19537\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__19534\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19531\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19522\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19519\
        );

    \I__1720\ : Span4Mux_h
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__1719\ : Span4Mux_s0_h
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__19513\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1717\ : InMux
    port map (
            O => \N__19510\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19504\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__19498\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19495\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1711\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19489\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__19483\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1707\ : InMux
    port map (
            O => \N__19480\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__19468\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1702\ : InMux
    port map (
            O => \N__19465\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19459\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__19456\,
            I => \N__19453\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__19453\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19436\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__19449\,
            I => \N__19433\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__19448\,
            I => \N__19430\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19427\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__19446\,
            I => \N__19424\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__19445\,
            I => \N__19421\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19418\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__19443\,
            I => \N__19415\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__19442\,
            I => \N__19412\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19409\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__19440\,
            I => \N__19406\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__19439\,
            I => \N__19403\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19400\
        );

    \I__1684\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19393\
        );

    \I__1683\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19393\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19393\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19384\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19384\
        );

    \I__1679\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19384\
        );

    \I__1678\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19384\
        );

    \I__1677\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19379\
        );

    \I__1676\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19379\
        );

    \I__1675\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19374\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19374\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__19400\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19393\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__19384\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__19379\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19374\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19363\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19360\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1666\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__19354\,
            I => un7_start_stop_0_a3
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19345\,
            I => \N__19342\
        );

    \I__1661\ : Span4Mux_h
    port map (
            O => \N__19342\,
            I => \N__19339\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__19339\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19336\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19330\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19327\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__19324\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__1653\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19315\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__19315\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19312\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19303\
        );

    \I__1648\ : Span4Mux_v
    port map (
            O => \N__19303\,
            I => \N__19300\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__19300\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19297\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1645\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__19288\,
            I => \N__19285\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__19285\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1641\ : InMux
    port map (
            O => \N__19282\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1640\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19276\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19276\,
            I => \N__19273\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__19273\,
            I => \N__19270\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__19270\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19267\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__19258\,
            I => \N__19255\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__19255\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1631\ : InMux
    port map (
            O => \N__19252\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1630\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19246\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__19246\,
            I => \N__19243\
        );

    \I__1628\ : Span4Mux_v
    port map (
            O => \N__19243\,
            I => \N__19240\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__19240\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1626\ : InMux
    port map (
            O => \N__19237\,
            I => \bfn_1_12_0_\
        );

    \I__1625\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19231\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19228\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__19225\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1621\ : InMux
    port map (
            O => \N__19222\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1620\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19216\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__19216\,
            I => \N__19213\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__19210\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1616\ : InMux
    port map (
            O => \N__19207\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1615\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__19195\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1611\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__19186\,
            I => \N__19183\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__19183\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__1606\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19174\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__19171\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19162\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__19159\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \N__19153\
        );

    \I__1598\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__19150\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1596\ : InMux
    port map (
            O => \N__19147\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1595\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19138\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__19138\,
            I => \N__19135\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__19135\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__1590\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19126\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__19126\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1588\ : InMux
    port map (
            O => \N__19123\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1587\ : IoInMux
    port map (
            O => \N__19120\,
            I => \N__19117\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__19117\,
            I => \N__19114\
        );

    \I__1585\ : Span4Mux_s3_v
    port map (
            O => \N__19114\,
            I => \N__19111\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__1583\ : Sp12to4
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__19102\,
            I => \N__19099\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__19099\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__1577\ : IoSpan4Mux
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__19084\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_16_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_27_0_\
        );

    \IN_MUX_bfv_16_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_16_28_0_\
        );

    \IN_MUX_bfv_16_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_16_29_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_13_27_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_17_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_17_27_0_\
        );

    \IN_MUX_bfv_17_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_17_28_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_12_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_26_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_8_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_8_24_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_7_17_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19120\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19096\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21124\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__46879\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__41269\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__40546\,
            CLKHFEN => \N__40612\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__40478\,
            RGB2PWM => \N__19957\,
            RGB1 => rgb_g_wire,
            CURREN => \N__40511\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19357\,
            RGB0PWM => \N__49555\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19204\,
            in2 => \_gnd_net_\,
            in3 => \N__19450\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19192\,
            in2 => \N__19180\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19168\,
            in2 => \N__19156\,
            in3 => \N__19147\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19144\,
            in2 => \N__19132\,
            in3 => \N__19123\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19333\,
            in2 => \N__19321\,
            in3 => \N__19312\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19309\,
            in2 => \N__19439\,
            in3 => \N__19297\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19294\,
            in2 => \N__19441\,
            in3 => \N__19282\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19279\,
            in2 => \N__19440\,
            in3 => \N__19267\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19264\,
            in2 => \N__19442\,
            in3 => \N__19252\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19249\,
            in2 => \N__19443\,
            in3 => \N__19237\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19234\,
            in2 => \N__19447\,
            in3 => \N__19222\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19219\,
            in2 => \N__19444\,
            in3 => \N__19207\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19507\,
            in2 => \N__19448\,
            in3 => \N__19495\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19492\,
            in2 => \N__19445\,
            in3 => \N__19480\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19477\,
            in2 => \N__19449\,
            in3 => \N__19465\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19462\,
            in2 => \N__19446\,
            in3 => \N__19363\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19360\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__43339\,
            in1 => \N__40317\,
            in2 => \_gnd_net_\,
            in3 => \N__42376\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_0_a3_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44812\,
            lcout => un7_start_stop_0_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39916\,
            in2 => \N__20235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37064\,
            in2 => \N__19351\,
            in3 => \N__19336\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37006\,
            in2 => \N__19681\,
            in3 => \N__19666\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36946\,
            in2 => \N__19663\,
            in3 => \N__19648\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36910\,
            in2 => \N__19645\,
            in3 => \N__19627\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36820\,
            in2 => \N__19624\,
            in3 => \N__19606\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37582\,
            in2 => \N__19603\,
            in3 => \N__19588\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37534\,
            in2 => \N__19585\,
            in3 => \N__19567\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37471\,
            in2 => \N__19564\,
            in3 => \N__19549\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37414\,
            in2 => \N__19546\,
            in3 => \N__19531\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37341\,
            in2 => \N__19528\,
            in3 => \N__19510\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37267\,
            in2 => \N__19813\,
            in3 => \N__19795\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37207\,
            in2 => \N__19792\,
            in3 => \N__19774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37153\,
            in2 => \N__19771\,
            in3 => \N__19753\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38029\,
            in2 => \N__19750\,
            in3 => \N__19735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19732\,
            in2 => \N__37983\,
            in3 => \N__19726\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19723\,
            in2 => \N__37926\,
            in3 => \N__19714\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37876\,
            in2 => \N__19711\,
            in3 => \N__19699\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37822\,
            in2 => \N__19696\,
            in3 => \N__19684\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37762\,
            in2 => \N__19948\,
            in3 => \N__19936\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37699\,
            in2 => \N__19933\,
            in3 => \N__19918\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37645\,
            in2 => \N__19915\,
            in3 => \N__19900\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38503\,
            in2 => \N__19897\,
            in3 => \N__19882\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38437\,
            in2 => \N__19879\,
            in3 => \N__19870\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38384\,
            in2 => \N__19867\,
            in3 => \N__19852\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38329\,
            in2 => \N__19849\,
            in3 => \N__19834\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38257\,
            in2 => \N__19831\,
            in3 => \N__19816\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38213\,
            in2 => \N__20068\,
            in3 => \N__20053\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38156\,
            in2 => \N__20050\,
            in3 => \N__20038\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38092\,
            in2 => \N__20035\,
            in3 => \N__20020\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20017\,
            in1 => \N__38708\,
            in2 => \N__20008\,
            in3 => \N__19993\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__20672\,
            in1 => \N__38730\,
            in2 => \N__19990\,
            in3 => \N__20377\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => 'H',
            sr => \N__49513\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011000101"
        )
    port map (
            in0 => \N__38729\,
            in1 => \N__19981\,
            in2 => \N__20426\,
            in3 => \N__20675\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => 'H',
            sr => \N__49513\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__38728\,
            in1 => \N__20674\,
            in2 => \N__20425\,
            in3 => \N__19972\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => 'H',
            sr => \N__49513\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__20673\,
            in1 => \N__38731\,
            in2 => \N__19966\,
            in3 => \N__20378\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49985\,
            ce => 'H',
            sr => \N__49513\
        );

    \phase_controller_inst1.N_39_i_i_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44811\,
            in2 => \_gnd_net_\,
            in3 => \N__49553\,
            lcout => \N_39_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20422\,
            in1 => \N__38803\,
            in2 => \N__20687\,
            in3 => \N__20134\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__20655\,
            in2 => \_gnd_net_\,
            in3 => \N__20423\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__38802\,
            in1 => \N__20656\,
            in2 => \N__20122\,
            in3 => \N__20424\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50013\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__20420\,
            in1 => \N__38779\,
            in2 => \N__20690\,
            in3 => \N__20113\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50005\,
            ce => 'H',
            sr => \N__49495\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__20419\,
            in1 => \_gnd_net_\,
            in2 => \N__20689\,
            in3 => \N__20104\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50005\,
            ce => 'H',
            sr => \N__49495\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__38777\,
            in1 => \N__20660\,
            in2 => \N__20098\,
            in3 => \N__20421\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50005\,
            ce => 'H',
            sr => \N__49495\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20418\,
            in1 => \N__38778\,
            in2 => \N__20688\,
            in3 => \N__20089\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50005\,
            ce => 'H',
            sr => \N__49495\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__38782\,
            in1 => \N__20403\,
            in2 => \N__20083\,
            in3 => \N__20652\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20650\,
            in1 => \N__38784\,
            in2 => \N__20434\,
            in3 => \N__20074\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__38783\,
            in1 => \N__20404\,
            in2 => \N__20203\,
            in3 => \N__20653\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001000"
        )
    port map (
            in0 => \N__20649\,
            in1 => \N__20194\,
            in2 => \N__20436\,
            in3 => \N__38786\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20651\,
            in1 => \N__38785\,
            in2 => \N__20435\,
            in3 => \N__20188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49996\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001000"
        )
    port map (
            in0 => \N__20398\,
            in1 => \N__20182\,
            in2 => \N__20691\,
            in3 => \N__38736\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__38733\,
            in1 => \N__20400\,
            in2 => \N__20176\,
            in3 => \N__20685\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20399\,
            in1 => \N__38735\,
            in2 => \N__20692\,
            in3 => \N__20167\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__38734\,
            in1 => \N__20401\,
            in2 => \N__20161\,
            in3 => \N__20686\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__38732\,
            in1 => \N__20678\,
            in2 => \N__20152\,
            in3 => \N__20402\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49986\,
            ce => 'H',
            sr => \N__49503\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20677\,
            in1 => \N__38738\,
            in2 => \N__20428\,
            in3 => \N__20140\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49509\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20676\,
            in1 => \N__38737\,
            in2 => \N__20427\,
            in3 => \N__20266\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49509\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38212\,
            in1 => \N__38383\,
            in2 => \N__38264\,
            in3 => \N__38333\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20260\,
            in1 => \N__20242\,
            in2 => \N__20254\,
            in3 => \N__20734\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37703\,
            in1 => \N__38699\,
            in2 => \N__38447\,
            in3 => \N__37763\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38040\,
            in1 => \N__37223\,
            in2 => \N__37427\,
            in3 => \N__37976\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38100\,
            in1 => \N__37287\,
            in2 => \N__20245\,
            in3 => \N__20275\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37925\,
            in1 => \N__37830\,
            in2 => \N__37656\,
            in3 => \N__37878\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37283\,
            in1 => \N__37340\,
            in2 => \N__37170\,
            in3 => \N__37975\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__20623\,
            in1 => \N__39915\,
            in2 => \N__20236\,
            in3 => \N__20433\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50006\,
            ce => 'H',
            sr => \N__49487\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20429\,
            in1 => \N__38792\,
            in2 => \N__20670\,
            in3 => \N__20212\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => 'H',
            sr => \N__49492\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__38790\,
            in1 => \N__20615\,
            in2 => \N__20515\,
            in3 => \N__20431\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => 'H',
            sr => \N__49492\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__20430\,
            in1 => \N__38793\,
            in2 => \N__20671\,
            in3 => \N__20503\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => 'H',
            sr => \N__49492\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__38791\,
            in1 => \N__20616\,
            in2 => \N__20494\,
            in3 => \N__20432\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49997\,
            ce => 'H',
            sr => \N__49492\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__20654\,
            in1 => \N__38781\,
            in2 => \N__20479\,
            in3 => \N__20417\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49987\,
            ce => 'H',
            sr => \N__49496\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20597\,
            in1 => \N__38799\,
            in2 => \N__20437\,
            in3 => \N__20464\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49974\,
            ce => 'H',
            sr => \N__49500\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__20598\,
            in2 => \N__20452\,
            in3 => \N__20385\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49963\,
            ce => 'H',
            sr => \N__49504\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37163\,
            in2 => \_gnd_net_\,
            in3 => \N__37330\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37536\,
            in1 => \N__37592\,
            in2 => \N__36848\,
            in3 => \N__37475\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__36965\,
            in1 => \N__37025\,
            in2 => \N__20269\,
            in3 => \N__36915\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38152\,
            in1 => \N__38504\,
            in2 => \N__20737\,
            in3 => \N__20728\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37924\,
            in1 => \N__37823\,
            in2 => \N__37655\,
            in3 => \N__37877\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38036\,
            in1 => \N__37224\,
            in2 => \N__37434\,
            in3 => \N__38157\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38337\,
            in2 => \_gnd_net_\,
            in3 => \N__37704\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__38448\,
            in1 => \N__37764\,
            in2 => \N__20722\,
            in3 => \N__20521\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__38511\,
            in1 => \N__38780\,
            in2 => \N__20719\,
            in3 => \N__20716\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20710\,
            in1 => \N__20701\,
            in2 => \N__20695\,
            in3 => \N__20767\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38220\,
            in1 => \N__38093\,
            in2 => \N__38271\,
            in3 => \N__38388\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26726\,
            in1 => \N__26707\,
            in2 => \_gnd_net_\,
            in3 => \N__30226\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50019\,
            ce => \N__29275\,
            sr => \N__49463\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27007\,
            in1 => \N__26963\,
            in2 => \_gnd_net_\,
            in3 => \N__30227\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50019\,
            ce => \N__29275\,
            sr => \N__49463\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30219\,
            in1 => \N__25994\,
            in2 => \_gnd_net_\,
            in3 => \N__26601\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__20794\,
            in1 => \N__25819\,
            in2 => \N__23164\,
            in3 => \N__27001\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26727\,
            in1 => \_gnd_net_\,
            in2 => \N__20755\,
            in3 => \N__26705\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20817\,
            in1 => \N__21565\,
            in2 => \_gnd_net_\,
            in3 => \N__30221\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30220\,
            in1 => \N__27002\,
            in2 => \_gnd_net_\,
            in3 => \N__26967\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__20778\,
            in1 => \N__23085\,
            in2 => \N__23119\,
            in3 => \N__20751\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__23118\,
            in1 => \N__20752\,
            in2 => \N__23086\,
            in3 => \N__20779\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30225\,
            in1 => \N__20813\,
            in2 => \_gnd_net_\,
            in3 => \N__21563\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50007\,
            ce => \N__29274\,
            sr => \N__49477\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27081\,
            in1 => \N__27053\,
            in2 => \_gnd_net_\,
            in3 => \N__30246\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49998\,
            ce => \N__29256\,
            sr => \N__49483\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30245\,
            in1 => \N__24900\,
            in2 => \_gnd_net_\,
            in3 => \N__24876\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49998\,
            ce => \N__29256\,
            sr => \N__49483\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27231\,
            in1 => \N__30247\,
            in2 => \_gnd_net_\,
            in3 => \N__27208\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49988\,
            ce => \N__29267\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26162\,
            in1 => \N__26141\,
            in2 => \_gnd_net_\,
            in3 => \N__30241\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24899\,
            in1 => \N__24875\,
            in2 => \_gnd_net_\,
            in3 => \N__30242\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27230\,
            in1 => \N__27206\,
            in2 => \_gnd_net_\,
            in3 => \N__30244\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27080\,
            in1 => \N__27057\,
            in2 => \_gnd_net_\,
            in3 => \N__30243\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__37035\,
            in1 => \N__37080\,
            in2 => \N__39942\,
            in3 => \N__36975\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__20761\,
            in1 => \N__37482\,
            in2 => \N__20770\,
            in3 => \N__36849\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__36914\,
            in1 => \N__37535\,
            in2 => \_gnd_net_\,
            in3 => \N__37593\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26914\,
            in1 => \N__26930\,
            in2 => \_gnd_net_\,
            in3 => \N__30319\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50014\,
            ce => \N__29235\,
            sr => \N__49438\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26068\,
            in1 => \N__26593\,
            in2 => \N__21564\,
            in3 => \N__26912\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30368\,
            in1 => \N__20821\,
            in2 => \_gnd_net_\,
            in3 => \N__21559\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50008\,
            ce => \N__30102\,
            sr => \N__49446\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26615\,
            in1 => \N__26519\,
            in2 => \N__28636\,
            in3 => \N__29494\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__24827\,
            in1 => \_gnd_net_\,
            in2 => \N__20797\,
            in3 => \N__30613\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21423\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49999\,
            ce => \N__22645\,
            sr => \N__49455\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21399\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49999\,
            ce => \N__22645\,
            sr => \N__49455\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26616\,
            in1 => \N__26645\,
            in2 => \_gnd_net_\,
            in3 => \N__30302\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22573\,
            in1 => \N__21419\,
            in2 => \_gnd_net_\,
            in3 => \N__20785\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22569\,
            in1 => \N__21395\,
            in2 => \_gnd_net_\,
            in3 => \N__20782\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22574\,
            in1 => \N__21376\,
            in2 => \_gnd_net_\,
            in3 => \N__20848\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22570\,
            in1 => \N__21354\,
            in2 => \_gnd_net_\,
            in3 => \N__20845\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22575\,
            in1 => \N__21332\,
            in2 => \_gnd_net_\,
            in3 => \N__20842\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22571\,
            in1 => \N__21306\,
            in2 => \_gnd_net_\,
            in3 => \N__20839\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22576\,
            in1 => \N__21286\,
            in2 => \_gnd_net_\,
            in3 => \N__20836\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22572\,
            in1 => \N__21268\,
            in2 => \_gnd_net_\,
            in3 => \N__20833\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__49989\,
            ce => \N__22410\,
            sr => \N__49464\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22564\,
            in1 => \N__21641\,
            in2 => \_gnd_net_\,
            in3 => \N__20830\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22568\,
            in1 => \N__21608\,
            in2 => \_gnd_net_\,
            in3 => \N__20827\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22561\,
            in1 => \N__21582\,
            in2 => \_gnd_net_\,
            in3 => \N__20824\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22565\,
            in1 => \N__21526\,
            in2 => \_gnd_net_\,
            in3 => \N__20875\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22562\,
            in1 => \N__21504\,
            in2 => \_gnd_net_\,
            in3 => \N__20872\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22566\,
            in1 => \N__21482\,
            in2 => \_gnd_net_\,
            in3 => \N__20869\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22563\,
            in1 => \N__21460\,
            in2 => \_gnd_net_\,
            in3 => \N__20866\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22567\,
            in1 => \N__21442\,
            in2 => \_gnd_net_\,
            in3 => \N__20863\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49975\,
            ce => \N__22411\,
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22529\,
            in1 => \N__21857\,
            in2 => \_gnd_net_\,
            in3 => \N__20860\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22548\,
            in1 => \N__21827\,
            in2 => \_gnd_net_\,
            in3 => \N__20857\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22530\,
            in1 => \N__21801\,
            in2 => \_gnd_net_\,
            in3 => \N__20854\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22549\,
            in1 => \N__21781\,
            in2 => \_gnd_net_\,
            in3 => \N__20851\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22531\,
            in1 => \N__21759\,
            in2 => \_gnd_net_\,
            in3 => \N__20902\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22550\,
            in1 => \N__21737\,
            in2 => \_gnd_net_\,
            in3 => \N__20899\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22532\,
            in1 => \N__21715\,
            in2 => \_gnd_net_\,
            in3 => \N__20896\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22551\,
            in1 => \N__21697\,
            in2 => \_gnd_net_\,
            in3 => \N__20893\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49964\,
            ce => \N__22409\,
            sr => \N__49478\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22542\,
            in1 => \N__21671\,
            in2 => \_gnd_net_\,
            in3 => \N__20890\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22546\,
            in1 => \N__21995\,
            in2 => \_gnd_net_\,
            in3 => \N__20887\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22543\,
            in1 => \N__21957\,
            in2 => \_gnd_net_\,
            in3 => \N__20884\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22547\,
            in1 => \N__21923\,
            in2 => \_gnd_net_\,
            in3 => \N__20881\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22544\,
            in1 => \N__21973\,
            in2 => \_gnd_net_\,
            in3 => \N__20878\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21937\,
            in1 => \N__22545\,
            in2 => \_gnd_net_\,
            in3 => \N__20932\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49955\,
            ce => \N__22399\,
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20929\,
            in2 => \_gnd_net_\,
            in3 => \N__21898\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21892\,
            in2 => \_gnd_net_\,
            in3 => \N__20923\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21883\,
            in2 => \_gnd_net_\,
            in3 => \N__20920\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21874\,
            in2 => \_gnd_net_\,
            in3 => \N__20917\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22078\,
            in2 => \_gnd_net_\,
            in3 => \N__20914\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22069\,
            in2 => \_gnd_net_\,
            in3 => \N__20911\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22060\,
            in2 => \_gnd_net_\,
            in3 => \N__20908\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22051\,
            in2 => \_gnd_net_\,
            in3 => \N__20905\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49489\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22042\,
            in2 => \_gnd_net_\,
            in3 => \N__20959\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22033\,
            in2 => \_gnd_net_\,
            in3 => \N__20956\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22024\,
            in2 => \_gnd_net_\,
            in3 => \N__20953\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22015\,
            in2 => \_gnd_net_\,
            in3 => \N__20950\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22006\,
            in2 => \_gnd_net_\,
            in3 => \N__20947\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22150\,
            in2 => \_gnd_net_\,
            in3 => \N__20944\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22141\,
            in2 => \_gnd_net_\,
            in3 => \N__20941\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22132\,
            in2 => \_gnd_net_\,
            in3 => \N__20938\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49493\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22123\,
            in2 => \_gnd_net_\,
            in3 => \N__20935\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22114\,
            in2 => \_gnd_net_\,
            in3 => \N__20986\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22105\,
            in2 => \_gnd_net_\,
            in3 => \N__20983\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22096\,
            in2 => \_gnd_net_\,
            in3 => \N__20980\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22087\,
            in2 => \_gnd_net_\,
            in3 => \N__20977\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22225\,
            in2 => \_gnd_net_\,
            in3 => \N__20974\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22216\,
            in2 => \_gnd_net_\,
            in3 => \N__20971\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22207\,
            in2 => \_gnd_net_\,
            in3 => \N__20968\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__49929\,
            ce => 'H',
            sr => \N__49497\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22198\,
            in2 => \_gnd_net_\,
            in3 => \N__20965\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22189\,
            in2 => \_gnd_net_\,
            in3 => \N__20962\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22180\,
            in2 => \_gnd_net_\,
            in3 => \N__21097\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22171\,
            in2 => \_gnd_net_\,
            in3 => \N__21094\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22162\,
            in2 => \_gnd_net_\,
            in3 => \N__21091\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22300\,
            in2 => \_gnd_net_\,
            in3 => \N__21088\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22255\,
            in2 => \_gnd_net_\,
            in3 => \N__21085\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22267\,
            in2 => \_gnd_net_\,
            in3 => \N__21082\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \N__49501\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21066\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49505\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21048\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49505\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => 'H',
            sr => \N__49510\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21006\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21186\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49514\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__22756\,
            in1 => \N__21144\,
            in2 => \_gnd_net_\,
            in3 => \N__21164\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21143\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__24054\,
            in1 => \N__42463\,
            in2 => \N__22762\,
            in3 => \N__21165\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.timer_s1.running_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__21166\,
            in1 => \N__22760\,
            in2 => \_gnd_net_\,
            in3 => \N__21145\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21163\,
            in2 => \_gnd_net_\,
            in3 => \N__21142\,
            lcout => \current_shift_inst.timer_s1.N_161_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22355\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => 'H',
            sr => \N__49415\
        );

    \delay_measurement_inst.stop_timer_hc_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22356\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => 'H',
            sr => \N__49415\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26072\,
            in1 => \N__26030\,
            in2 => \_gnd_net_\,
            in3 => \N__30330\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__23061\,
            in1 => \N__21250\,
            in2 => \N__23035\,
            in3 => \N__21235\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30329\,
            in1 => \N__26934\,
            in2 => \_gnd_net_\,
            in3 => \N__26911\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__21249\,
            in1 => \N__23028\,
            in2 => \N__23062\,
            in3 => \N__21234\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26860\,
            in1 => \N__26820\,
            in2 => \_gnd_net_\,
            in3 => \N__30303\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => \elapsed_time_ns_1_RNI46CN9_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30304\,
            in1 => \_gnd_net_\,
            in2 => \N__21238\,
            in3 => \N__26861\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50009\,
            ce => \N__29215\,
            sr => \N__49430\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26001\,
            in1 => \N__26594\,
            in2 => \_gnd_net_\,
            in3 => \N__30305\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50009\,
            ce => \N__29215\,
            sr => \N__49430\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__21220\,
            in1 => \N__22983\,
            in2 => \N__21211\,
            in3 => \N__23001\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26792\,
            in1 => \N__26754\,
            in2 => \_gnd_net_\,
            in3 => \N__30356\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30357\,
            in1 => \_gnd_net_\,
            in2 => \N__21223\,
            in3 => \N__26793\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50000\,
            ce => \N__29255\,
            sr => \N__49439\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__21219\,
            in1 => \N__22982\,
            in2 => \N__21210\,
            in3 => \N__23000\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21374\,
            in2 => \N__21424\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21353\,
            in2 => \N__21403\,
            in3 => \N__21379\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21375\,
            in2 => \N__21333\,
            in3 => \N__21361\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21305\,
            in2 => \N__21358\,
            in3 => \N__21337\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21284\,
            in2 => \N__21334\,
            in3 => \N__21313\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21266\,
            in2 => \N__21310\,
            in3 => \N__21289\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21285\,
            in2 => \N__21649\,
            in3 => \N__21271\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21267\,
            in2 => \N__21619\,
            in3 => \N__21253\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49990\,
            ce => \N__22644\,
            sr => \N__49447\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21581\,
            in2 => \N__21648\,
            in3 => \N__21622\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21524\,
            in2 => \N__21615\,
            in3 => \N__21589\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21503\,
            in2 => \N__21586\,
            in3 => \N__21529\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21525\,
            in2 => \N__21483\,
            in3 => \N__21511\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21458\,
            in2 => \N__21508\,
            in3 => \N__21487\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21440\,
            in2 => \N__21484\,
            in3 => \N__21463\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21459\,
            in2 => \N__21865\,
            in3 => \N__21445\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21441\,
            in2 => \N__21835\,
            in3 => \N__21427\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49976\,
            ce => \N__22643\,
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21800\,
            in2 => \N__21864\,
            in3 => \N__21838\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21779\,
            in2 => \N__21834\,
            in3 => \N__21808\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21758\,
            in2 => \N__21805\,
            in3 => \N__21784\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21780\,
            in2 => \N__21738\,
            in3 => \N__21766\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21713\,
            in2 => \N__21763\,
            in3 => \N__21742\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21695\,
            in2 => \N__21739\,
            in3 => \N__21718\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21714\,
            in2 => \N__21679\,
            in3 => \N__21700\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21696\,
            in2 => \N__22000\,
            in3 => \N__21682\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49965\,
            ce => \N__22642\,
            sr => \N__49465\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21956\,
            in2 => \N__21678\,
            in3 => \N__21652\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49956\,
            ce => \N__22629\,
            sr => \N__49470\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21996\,
            in2 => \N__21924\,
            in3 => \N__21976\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49956\,
            ce => \N__22629\,
            sr => \N__49470\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21972\,
            in2 => \N__21961\,
            in3 => \N__21940\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49956\,
            ce => \N__22629\,
            sr => \N__49470\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21936\,
            in2 => \N__21925\,
            in3 => \N__21904\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49956\,
            ce => \N__22629\,
            sr => \N__49470\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21901\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__22629\,
            sr => \N__49470\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23302\,
            in2 => \N__23290\,
            in3 => \N__23288\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23380\,
            in2 => \_gnd_net_\,
            in3 => \N__21886\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23251\,
            in2 => \_gnd_net_\,
            in3 => \N__21877\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23257\,
            in2 => \_gnd_net_\,
            in3 => \N__21868\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23368\,
            in2 => \_gnd_net_\,
            in3 => \N__22072\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23362\,
            in2 => \_gnd_net_\,
            in3 => \N__22063\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23356\,
            in2 => \_gnd_net_\,
            in3 => \N__22054\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22423\,
            in2 => \_gnd_net_\,
            in3 => \N__22045\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23320\,
            in2 => \_gnd_net_\,
            in3 => \N__22036\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23269\,
            in2 => \_gnd_net_\,
            in3 => \N__22027\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23350\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23263\,
            in2 => \_gnd_net_\,
            in3 => \N__22009\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23338\,
            in2 => \_gnd_net_\,
            in3 => \N__22153\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23344\,
            in2 => \_gnd_net_\,
            in3 => \N__22144\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23326\,
            in2 => \_gnd_net_\,
            in3 => \N__22135\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23404\,
            in2 => \_gnd_net_\,
            in3 => \N__22126\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23374\,
            in2 => \_gnd_net_\,
            in3 => \N__22117\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22441\,
            in2 => \_gnd_net_\,
            in3 => \N__22108\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22288\,
            in2 => \_gnd_net_\,
            in3 => \N__22099\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22432\,
            in2 => \_gnd_net_\,
            in3 => \N__22090\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23332\,
            in2 => \_gnd_net_\,
            in3 => \N__22081\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22276\,
            in2 => \_gnd_net_\,
            in3 => \N__22219\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22249\,
            in2 => \_gnd_net_\,
            in3 => \N__22210\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22240\,
            in2 => \_gnd_net_\,
            in3 => \N__22201\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22231\,
            in2 => \_gnd_net_\,
            in3 => \N__22192\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22582\,
            in2 => \_gnd_net_\,
            in3 => \N__22183\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23398\,
            in3 => \N__22174\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22282\,
            in2 => \_gnd_net_\,
            in3 => \N__22165\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25243\,
            in2 => \_gnd_net_\,
            in3 => \N__22156\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23314\,
            in2 => \_gnd_net_\,
            in3 => \N__22294\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \_gnd_net_\,
            in3 => \N__22291\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__25376\,
            in1 => \N__25009\,
            in2 => \_gnd_net_\,
            in3 => \N__27988\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25352\,
            in1 => \N__28090\,
            in2 => \_gnd_net_\,
            in3 => \N__25390\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27928\,
            in1 => \N__25156\,
            in2 => \_gnd_net_\,
            in3 => \N__25347\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__27913\,
            in2 => \_gnd_net_\,
            in3 => \N__25144\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25132\,
            in1 => \N__27883\,
            in2 => \_gnd_net_\,
            in3 => \N__25349\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25350\,
            in1 => \N__28138\,
            in2 => \_gnd_net_\,
            in3 => \N__25120\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__25108\,
            in1 => \N__25351\,
            in2 => \_gnd_net_\,
            in3 => \N__28123\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__28003\,
            in1 => \N__25024\,
            in2 => \_gnd_net_\,
            in3 => \N__25294\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__25295\,
            in1 => \N__25180\,
            in2 => \_gnd_net_\,
            in3 => \N__27958\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35551\,
            in1 => \N__25758\,
            in2 => \N__35237\,
            in3 => \N__28459\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32778\,
            in1 => \N__31952\,
            in2 => \_gnd_net_\,
            in3 => \N__31989\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27595\,
            in1 => \N__24949\,
            in2 => \_gnd_net_\,
            in3 => \N__25293\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__22334\,
            in2 => \_gnd_net_\,
            in3 => \N__22362\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__22363\,
            in1 => \_gnd_net_\,
            in2 => \N__22339\,
            in3 => \N__22318\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49506\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22316\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__48554\,
            in2 => \_gnd_net_\,
            in3 => \N__48516\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32248\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35602\,
            in2 => \N__22597\,
            in3 => \N__32953\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32183\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__32881\,
            sr => \N__49511\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32211\,
            in1 => \N__40616\,
            in2 => \_gnd_net_\,
            in3 => \N__22594\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__40617\,
            in1 => \_gnd_net_\,
            in2 => \N__22588\,
            in3 => \N__27501\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32489\,
            in1 => \N__32777\,
            in2 => \_gnd_net_\,
            in3 => \N__32469\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32488\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22921\,
            in1 => \N__32970\,
            in2 => \_gnd_net_\,
            in3 => \N__22585\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22917\,
            in1 => \N__32898\,
            in2 => \_gnd_net_\,
            in3 => \N__22672\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_2_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22922\,
            in1 => \N__23618\,
            in2 => \_gnd_net_\,
            in3 => \N__22669\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_3_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22918\,
            in1 => \N__23588\,
            in2 => \_gnd_net_\,
            in3 => \N__22666\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_4_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22923\,
            in1 => \N__23568\,
            in2 => \_gnd_net_\,
            in3 => \N__22663\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_5_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22919\,
            in1 => \N__23544\,
            in2 => \_gnd_net_\,
            in3 => \N__22660\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_6_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22924\,
            in1 => \N__23521\,
            in2 => \_gnd_net_\,
            in3 => \N__22657\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_7_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22920\,
            in1 => \N__23503\,
            in2 => \_gnd_net_\,
            in3 => \N__22654\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49894\,
            ce => \N__22798\,
            sr => \N__49515\
        );

    \current_shift_inst.timer_s1.counter_8_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22912\,
            in1 => \N__23477\,
            in2 => \_gnd_net_\,
            in3 => \N__22651\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_9_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22916\,
            in1 => \N__23447\,
            in2 => \_gnd_net_\,
            in3 => \N__22648\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_10_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22909\,
            in1 => \N__23832\,
            in2 => \_gnd_net_\,
            in3 => \N__22699\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_11_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22913\,
            in1 => \N__23809\,
            in2 => \_gnd_net_\,
            in3 => \N__22696\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_12_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22910\,
            in1 => \N__23790\,
            in2 => \_gnd_net_\,
            in3 => \N__22693\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_13_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22914\,
            in1 => \N__23765\,
            in2 => \_gnd_net_\,
            in3 => \N__22690\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_14_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22911\,
            in1 => \N__23743\,
            in2 => \_gnd_net_\,
            in3 => \N__22687\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_15_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22915\,
            in1 => \N__23725\,
            in2 => \_gnd_net_\,
            in3 => \N__22684\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49887\,
            ce => \N__22797\,
            sr => \N__49519\
        );

    \current_shift_inst.timer_s1.counter_16_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22881\,
            in1 => \N__23702\,
            in2 => \_gnd_net_\,
            in3 => \N__22681\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_17_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22885\,
            in1 => \N__23669\,
            in2 => \_gnd_net_\,
            in3 => \N__22678\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_18_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22882\,
            in1 => \N__23643\,
            in2 => \_gnd_net_\,
            in3 => \N__22675\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_19_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22886\,
            in1 => \N__24031\,
            in2 => \_gnd_net_\,
            in3 => \N__22726\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_20_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22883\,
            in1 => \N__24012\,
            in2 => \_gnd_net_\,
            in3 => \N__22723\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_21_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22887\,
            in1 => \N__23987\,
            in2 => \_gnd_net_\,
            in3 => \N__22720\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_22_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22884\,
            in1 => \N__23965\,
            in2 => \_gnd_net_\,
            in3 => \N__22717\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_23_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22888\,
            in1 => \N__23947\,
            in2 => \_gnd_net_\,
            in3 => \N__22714\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49882\,
            ce => \N__22784\,
            sr => \N__49522\
        );

    \current_shift_inst.timer_s1.counter_24_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22877\,
            in1 => \N__23924\,
            in2 => \_gnd_net_\,
            in3 => \N__22711\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.timer_s1.counter_25_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22889\,
            in1 => \N__23894\,
            in2 => \_gnd_net_\,
            in3 => \N__22708\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.timer_s1.counter_26_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22878\,
            in1 => \N__23856\,
            in2 => \_gnd_net_\,
            in3 => \N__22705\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.timer_s1.counter_27_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22890\,
            in1 => \N__24090\,
            in2 => \_gnd_net_\,
            in3 => \N__22702\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.timer_s1.counter_28_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22879\,
            in1 => \N__23869\,
            in2 => \_gnd_net_\,
            in3 => \N__22927\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.timer_s1.counter_29_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24103\,
            in1 => \N__22880\,
            in2 => \_gnd_net_\,
            in3 => \N__22801\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => \N__22783\,
            sr => \N__49524\
        );

    \current_shift_inst.start_timer_s1_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__22761\,
            in2 => \_gnd_net_\,
            in3 => \N__42461\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => 'H',
            sr => \N__49526\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26452\,
            in1 => \N__26409\,
            in2 => \_gnd_net_\,
            in3 => \N__30328\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24193\,
            in2 => \N__25849\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29186\,
            in1 => \N__24172\,
            in2 => \_gnd_net_\,
            in3 => \N__22738\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29190\,
            in1 => \N__24151\,
            in2 => \N__24205\,
            in3 => \N__22735\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29187\,
            in1 => \N__24124\,
            in2 => \_gnd_net_\,
            in3 => \N__22732\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29191\,
            in1 => \N__24370\,
            in2 => \_gnd_net_\,
            in3 => \N__22729\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29188\,
            in1 => \N__24349\,
            in2 => \_gnd_net_\,
            in3 => \N__22954\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29192\,
            in1 => \N__24331\,
            in2 => \_gnd_net_\,
            in3 => \N__22951\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29189\,
            in1 => \N__24310\,
            in2 => \_gnd_net_\,
            in3 => \N__22948\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__50001\,
            ce => 'H',
            sr => \N__49423\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29124\,
            in1 => \N__24292\,
            in2 => \_gnd_net_\,
            in3 => \N__22945\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29117\,
            in1 => \N__24274\,
            in2 => \_gnd_net_\,
            in3 => \N__22942\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29121\,
            in1 => \N__24256\,
            in2 => \_gnd_net_\,
            in3 => \N__22939\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29118\,
            in1 => \N__24232\,
            in2 => \_gnd_net_\,
            in3 => \N__22936\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29122\,
            in1 => \N__24538\,
            in2 => \_gnd_net_\,
            in3 => \N__22933\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29119\,
            in1 => \N__24502\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29123\,
            in1 => \N__24472\,
            in2 => \_gnd_net_\,
            in3 => \N__23065\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29120\,
            in1 => \N__23060\,
            in2 => \_gnd_net_\,
            in3 => \N__23038\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49991\,
            ce => 'H',
            sr => \N__49431\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29193\,
            in1 => \N__23027\,
            in2 => \_gnd_net_\,
            in3 => \N__23005\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29239\,
            in1 => \N__23002\,
            in2 => \_gnd_net_\,
            in3 => \N__22987\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29194\,
            in1 => \N__22984\,
            in2 => \_gnd_net_\,
            in3 => \N__22969\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29240\,
            in1 => \N__25931\,
            in2 => \_gnd_net_\,
            in3 => \N__22966\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29195\,
            in1 => \N__25952\,
            in2 => \_gnd_net_\,
            in3 => \N__22963\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29241\,
            in1 => \N__24692\,
            in2 => \_gnd_net_\,
            in3 => \N__22960\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29196\,
            in1 => \N__24710\,
            in2 => \_gnd_net_\,
            in3 => \N__22957\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29242\,
            in1 => \N__23195\,
            in2 => \_gnd_net_\,
            in3 => \N__23137\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29223\,
            in1 => \N__23233\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29236\,
            in1 => \N__24574\,
            in2 => \_gnd_net_\,
            in3 => \N__23131\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29224\,
            in1 => \N__24591\,
            in2 => \_gnd_net_\,
            in3 => \N__23128\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29237\,
            in1 => \N__26210\,
            in2 => \_gnd_net_\,
            in3 => \N__23125\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29225\,
            in1 => \N__26231\,
            in2 => \_gnd_net_\,
            in3 => \N__23122\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29238\,
            in1 => \N__23108\,
            in2 => \_gnd_net_\,
            in3 => \N__23092\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29226\,
            in1 => \N__23081\,
            in2 => \_gnd_net_\,
            in3 => \N__23089\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49966\,
            ce => 'H',
            sr => \N__49448\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__23242\,
            in1 => \N__23232\,
            in2 => \N__23218\,
            in3 => \N__23197\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26321\,
            in1 => \N__26298\,
            in2 => \_gnd_net_\,
            in3 => \N__30526\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30527\,
            in1 => \_gnd_net_\,
            in2 => \N__23245\,
            in3 => \N__26322\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49957\,
            ce => \N__29266\,
            sr => \N__49457\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__23241\,
            in1 => \N__23231\,
            in2 => \N__23217\,
            in3 => \N__23196\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26791\,
            in1 => \N__26686\,
            in2 => \N__26865\,
            in3 => \N__29447\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23149\,
            in1 => \N__23143\,
            in2 => \N__23179\,
            in3 => \N__23176\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28995\,
            in2 => \N__48571\,
            in3 => \N__48517\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__24856\,
            in2 => \N__26131\,
            in3 => \N__27040\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26380\,
            in1 => \N__26342\,
            in2 => \_gnd_net_\,
            in3 => \N__30346\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27187\,
            in1 => \N__27267\,
            in2 => \N__26480\,
            in3 => \N__26320\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24934\,
            in1 => \N__27868\,
            in2 => \_gnd_net_\,
            in3 => \N__25358\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24790\,
            in1 => \N__27721\,
            in2 => \_gnd_net_\,
            in3 => \N__25356\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23293\,
            in3 => \N__23289\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49471\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25357\,
            lcout => \current_shift_inst.N_1306_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25359\,
            in1 => \N__27850\,
            in2 => \_gnd_net_\,
            in3 => \N__24922\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__25367\,
            in1 => \N__25081\,
            in2 => \_gnd_net_\,
            in3 => \N__27811\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__24988\,
            in1 => \N__25363\,
            in2 => \_gnd_net_\,
            in3 => \N__27667\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25362\,
            in1 => \N__27682\,
            in2 => \_gnd_net_\,
            in3 => \N__24997\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27703\,
            in1 => \N__24781\,
            in2 => \_gnd_net_\,
            in3 => \N__25361\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25368\,
            in1 => \N__28030\,
            in2 => \_gnd_net_\,
            in3 => \N__25036\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27652\,
            in1 => \N__24976\,
            in2 => \_gnd_net_\,
            in3 => \N__25364\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__24967\,
            in2 => \_gnd_net_\,
            in3 => \N__27634\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27616\,
            in1 => \N__24958\,
            in2 => \_gnd_net_\,
            in3 => \N__25366\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__24910\,
            in1 => \N__27826\,
            in2 => \_gnd_net_\,
            in3 => \N__25369\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__25371\,
            in1 => \N__25063\,
            in2 => \_gnd_net_\,
            in3 => \N__27778\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27796\,
            in1 => \N__25072\,
            in2 => \_gnd_net_\,
            in3 => \N__25370\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25374\,
            in1 => \N__27943\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27760\,
            in1 => \N__25054\,
            in2 => \_gnd_net_\,
            in3 => \N__25372\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__25373\,
            in1 => \N__27739\,
            in2 => \_gnd_net_\,
            in3 => \N__25045\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__28108\,
            in1 => \N__25093\,
            in2 => \_gnd_net_\,
            in3 => \N__25375\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32584\,
            in2 => \N__32215\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40732\,
            in2 => \N__32617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25549\,
            in2 => \N__40755\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40736\,
            in2 => \N__25486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25561\,
            in2 => \N__40756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40740\,
            in2 => \N__27448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23389\,
            in2 => \N__40757\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40744\,
            in2 => \N__27427\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40728\,
            in2 => \N__31834\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32263\,
            in2 => \N__40754\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40716\,
            in2 => \N__25198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23416\,
            in2 => \N__40751\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40720\,
            in2 => \N__25471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25222\,
            in2 => \N__40752\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40724\,
            in2 => \N__25216\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25588\,
            in2 => \N__40753\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40659\,
            in2 => \N__25462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25231\,
            in2 => \N__40712\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40663\,
            in2 => \N__25663\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25414\,
            in2 => \N__40713\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40667\,
            in2 => \N__25645\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25789\,
            in2 => \N__40714\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40671\,
            in2 => \N__25408\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25189\,
            in2 => \N__40715\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40618\,
            in2 => \N__25576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25537\,
            in2 => \N__40656\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40622\,
            in2 => \N__25681\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25435\,
            in2 => \N__40657\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40626\,
            in2 => \N__25453\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25516\,
            in2 => \N__40658\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40630\,
            in2 => \N__25444\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35595\,
            in2 => \_gnd_net_\,
            in3 => \N__23422\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32969\,
            in2 => \N__23619\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32897\,
            in2 => \N__23595\,
            in3 => \N__23419\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \N__23620\,
            in3 => \N__23599\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23540\,
            in2 => \N__23596\,
            in3 => \N__23572\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23519\,
            in2 => \N__23569\,
            in3 => \N__23548\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23501\,
            in2 => \N__23545\,
            in3 => \N__23524\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23520\,
            in2 => \N__23485\,
            in3 => \N__23506\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23502\,
            in2 => \N__23452\,
            in3 => \N__23488\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49895\,
            ce => \N__32880\,
            sr => \N__49507\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23828\,
            in2 => \N__23481\,
            in3 => \N__23455\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23807\,
            in2 => \N__23451\,
            in3 => \N__23425\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23786\,
            in2 => \N__23833\,
            in3 => \N__23812\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23808\,
            in2 => \N__23766\,
            in3 => \N__23794\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23741\,
            in2 => \N__23791\,
            in3 => \N__23770\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23723\,
            in2 => \N__23767\,
            in3 => \N__23746\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23742\,
            in2 => \N__23707\,
            in3 => \N__23728\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23724\,
            in2 => \N__23676\,
            in3 => \N__23710\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49888\,
            ce => \N__32879\,
            sr => \N__49512\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23639\,
            in2 => \N__23706\,
            in3 => \N__23680\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24029\,
            in2 => \N__23677\,
            in3 => \N__23647\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24008\,
            in2 => \N__23644\,
            in3 => \N__23623\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24030\,
            in2 => \N__23988\,
            in3 => \N__24016\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23963\,
            in2 => \N__24013\,
            in3 => \N__23992\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23945\,
            in2 => \N__23989\,
            in3 => \N__23968\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23964\,
            in2 => \N__23929\,
            in3 => \N__23950\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23946\,
            in2 => \N__23899\,
            in3 => \N__23932\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49883\,
            ce => \N__32877\,
            sr => \N__49516\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23852\,
            in2 => \N__23928\,
            in3 => \N__23902\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49879\,
            ce => \N__32876\,
            sr => \N__49520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24086\,
            in2 => \N__23898\,
            in3 => \N__23872\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49879\,
            ce => \N__32876\,
            sr => \N__49520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23868\,
            in2 => \N__23857\,
            in3 => \N__23836\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49879\,
            ce => \N__32876\,
            sr => \N__49520\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24102\,
            in2 => \N__24091\,
            in3 => \N__24070\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49879\,
            ce => \N__32876\,
            sr => \N__49520\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24067\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31348\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42462\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => 'H',
            sr => \N__49525\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28668\,
            in1 => \N__28650\,
            in2 => \_gnd_net_\,
            in3 => \N__30432\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50002\,
            ce => \N__29219\,
            sr => \N__49397\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30421\,
            in1 => \N__26555\,
            in2 => \_gnd_net_\,
            in3 => \N__26538\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49992\,
            ce => \N__29246\,
            sr => \N__49403\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26460\,
            in1 => \N__26405\,
            in2 => \_gnd_net_\,
            in3 => \N__30423\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49992\,
            ce => \N__29246\,
            sr => \N__49403\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26034\,
            in1 => \N__26076\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49992\,
            ce => \N__29246\,
            sr => \N__49403\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28994\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__37125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28577\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__28575\,
            in1 => \N__25872\,
            in2 => \_gnd_net_\,
            in3 => \N__37124\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24208\,
            in3 => \N__25860\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__28576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28547\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24196\,
            in3 => \N__28603\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24187\,
            in2 => \N__25882\,
            in3 => \N__25838\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24181\,
            in2 => \N__24160\,
            in3 => \N__24171\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24139\,
            in2 => \N__24655\,
            in3 => \N__24150\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24133\,
            in2 => \N__24112\,
            in3 => \N__24123\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24379\,
            in2 => \N__24358\,
            in3 => \N__24369\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24337\,
            in2 => \N__24604\,
            in3 => \N__24348\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26185\,
            in2 => \N__24319\,
            in3 => \N__24330\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24298\,
            in2 => \N__29290\,
            in3 => \N__24309\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24291\,
            in1 => \N__24280\,
            in2 => \N__25978\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24262\,
            in2 => \N__25798\,
            in3 => \N__24273\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25969\,
            in2 => \N__24244\,
            in3 => \N__24255\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29299\,
            in2 => \N__24220\,
            in3 => \N__24231\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24553\,
            in2 => \N__24526\,
            in3 => \N__24537\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24514\,
            in2 => \N__24490\,
            in3 => \N__24501\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24481\,
            in2 => \N__24460\,
            in3 => \N__24471\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24451\,
            in2 => \N__24439\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24424\,
            in2 => \N__24412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25915\,
            in2 => \N__25963\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24676\,
            in2 => \N__24745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24397\,
            in2 => \N__24388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24559\,
            in2 => \N__24616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26194\,
            in2 => \N__26245\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24643\,
            in2 => \N__24631\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24619\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__24573\,
            in1 => \N__24754\,
            in2 => \N__24769\,
            in3 => \N__24590\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30501\,
            in1 => \N__26285\,
            in2 => \_gnd_net_\,
            in3 => \N__26256\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26286\,
            in1 => \_gnd_net_\,
            in2 => \N__24607\,
            in3 => \N__30504\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49942\,
            ce => \N__29265\,
            sr => \N__49441\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__24753\,
            in1 => \N__24768\,
            in2 => \N__24592\,
            in3 => \N__24572\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24836\,
            in1 => \N__24801\,
            in2 => \_gnd_net_\,
            in3 => \N__30500\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30503\,
            in1 => \_gnd_net_\,
            in2 => \N__24772\,
            in3 => \N__24837\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49942\,
            ce => \N__29265\,
            sr => \N__49441\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30668\,
            in1 => \N__30639\,
            in2 => \_gnd_net_\,
            in3 => \N__30499\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30502\,
            in1 => \_gnd_net_\,
            in2 => \N__24757\,
            in3 => \N__30669\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49942\,
            ce => \N__29265\,
            sr => \N__49441\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__24694\,
            in1 => \N__24664\,
            in2 => \N__24730\,
            in3 => \N__24714\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__24663\,
            in1 => \N__24729\,
            in2 => \N__24715\,
            in3 => \N__24693\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27281\,
            in1 => \N__27252\,
            in2 => \_gnd_net_\,
            in3 => \N__30429\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30430\,
            in1 => \_gnd_net_\,
            in2 => \N__24667\,
            in3 => \N__27282\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49931\,
            ce => \N__29254\,
            sr => \N__49449\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26652\,
            in1 => \N__26628\,
            in2 => \_gnd_net_\,
            in3 => \N__30431\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49931\,
            ce => \N__29254\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30426\,
            in1 => \N__26169\,
            in2 => \_gnd_net_\,
            in3 => \N__26143\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__30097\,
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27116\,
            in1 => \_gnd_net_\,
            in2 => \N__27157\,
            in3 => \N__30427\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__30097\,
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24901\,
            in1 => \N__24877\,
            in2 => \_gnd_net_\,
            in3 => \N__30428\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__30097\,
            sr => \N__49458\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30425\,
            in1 => \N__24838\,
            in2 => \_gnd_net_\,
            in3 => \N__24805\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__30097\,
            sr => \N__49458\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25498\,
            in2 => \N__27535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32822\,
            in2 => \N__32926\,
            in3 => \N__32596\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32597\,
            in1 => \N__34719\,
            in2 => \N__30931\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31000\,
            in2 => \N__34869\,
            in3 => \N__24784\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34723\,
            in2 => \N__25531\,
            in3 => \N__24775\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25399\,
            in2 => \N__34870\,
            in3 => \N__24991\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34727\,
            in2 => \N__25429\,
            in3 => \N__24979\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31744\,
            in2 => \N__34871\,
            in3 => \N__24970\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34731\,
            in2 => \N__27487\,
            in3 => \N__24961\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32347\,
            in2 => \N__34872\,
            in3 => \N__24952\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34735\,
            in2 => \N__27547\,
            in3 => \N__24937\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25600\,
            in2 => \N__34873\,
            in3 => \N__24925\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34739\,
            in2 => \N__27436\,
            in3 => \N__24913\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25609\,
            in2 => \N__34874\,
            in3 => \N__24904\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34743\,
            in2 => \N__27358\,
            in3 => \N__25075\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26947\,
            in2 => \N__34875\,
            in3 => \N__25066\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34977\,
            in2 => \N__27295\,
            in3 => \N__25057\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27577\,
            in2 => \N__35136\,
            in3 => \N__25048\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34981\,
            in2 => \N__25696\,
            in3 => \N__25039\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27583\,
            in2 => \N__35137\,
            in3 => \N__25027\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34985\,
            in2 => \N__27304\,
            in3 => \N__25012\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27346\,
            in2 => \N__35138\,
            in3 => \N__25000\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34989\,
            in2 => \N__27367\,
            in3 => \N__25168\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27571\,
            in2 => \N__35139\,
            in3 => \N__25159\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35000\,
            in2 => \N__27565\,
            in3 => \N__25147\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25777\,
            in2 => \N__35143\,
            in3 => \N__25135\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35004\,
            in2 => \N__25729\,
            in3 => \N__25123\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27556\,
            in2 => \N__35144\,
            in3 => \N__25111\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35008\,
            in2 => \N__25714\,
            in3 => \N__25096\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25768\,
            in2 => \N__35145\,
            in3 => \N__25084\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35012\,
            in2 => \N__25207\,
            in3 => \N__25381\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__32320\,
            in1 => \N__28069\,
            in2 => \N__25378\,
            in3 => \N__25246\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32783\,
            in1 => \N__31358\,
            in2 => \_gnd_net_\,
            in3 => \N__31401\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__25630\,
            in1 => \N__35534\,
            in2 => \N__28387\,
            in3 => \N__35184\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32781\,
            in1 => \N__25629\,
            in2 => \_gnd_net_\,
            in3 => \N__28383\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31079\,
            in1 => \N__32782\,
            in2 => \_gnd_net_\,
            in3 => \N__30908\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__35185\,
            in1 => \N__35535\,
            in2 => \N__32598\,
            in3 => \N__32542\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32138\,
            in1 => \N__32779\,
            in2 => \_gnd_net_\,
            in3 => \N__32113\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__32784\,
            in1 => \N__34637\,
            in2 => \_gnd_net_\,
            in3 => \N__35283\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__31684\,
            in1 => \N__32780\,
            in2 => \_gnd_net_\,
            in3 => \N__31715\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32761\,
            in1 => \N__30854\,
            in2 => \_gnd_net_\,
            in3 => \N__30809\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31302\,
            in1 => \N__35574\,
            in2 => \_gnd_net_\,
            in3 => \N__31269\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35576\,
            in1 => \N__35148\,
            in2 => \N__28254\,
            in3 => \N__27474\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32541\,
            in2 => \_gnd_net_\,
            in3 => \N__35575\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35573\,
            in1 => \N__28856\,
            in2 => \_gnd_net_\,
            in3 => \N__28818\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35149\,
            in1 => \N__35577\,
            in2 => \N__31956\,
            in3 => \N__31985\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32762\,
            in1 => \N__31628\,
            in2 => \_gnd_net_\,
            in3 => \N__31599\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27411\,
            in1 => \N__32763\,
            in2 => \_gnd_net_\,
            in3 => \N__28518\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__27473\,
            in1 => \N__35580\,
            in2 => \N__28255\,
            in3 => \N__35076\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35552\,
            in1 => \N__31523\,
            in2 => \_gnd_net_\,
            in3 => \N__31557\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35579\,
            in1 => \N__31222\,
            in2 => \N__35192\,
            in3 => \N__31200\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32286\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35578\,
            in1 => \N__28770\,
            in2 => \_gnd_net_\,
            in3 => \N__28741\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31760\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__25507\,
            in1 => \N__35553\,
            in2 => \_gnd_net_\,
            in3 => \N__32952\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__28299\,
            in1 => \N__35583\,
            in2 => \N__35193\,
            in3 => \N__27329\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32743\,
            in1 => \N__30972\,
            in2 => \_gnd_net_\,
            in3 => \N__30948\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27469\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30971\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31942\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31457\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__31227\,
            in1 => \N__32744\,
            in2 => \N__31199\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31226\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32708\,
            in1 => \N__31475\,
            in2 => \_gnd_net_\,
            in3 => \N__31430\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32129\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31705\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25622\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__25623\,
            in1 => \N__35582\,
            in2 => \N__28382\,
            in3 => \N__35197\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35581\,
            in1 => \N__32490\,
            in2 => \N__35238\,
            in3 => \N__32462\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32709\,
            in1 => \N__31142\,
            in2 => \_gnd_net_\,
            in3 => \N__31103\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31141\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32369\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32788\,
            in1 => \N__32023\,
            in2 => \_gnd_net_\,
            in3 => \N__32052\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27385\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30751\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31619\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27322\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35266\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30844\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35198\,
            in1 => \N__35604\,
            in2 => \N__30768\,
            in3 => \N__30729\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35603\,
            in1 => \N__25745\,
            in2 => \_gnd_net_\,
            in3 => \N__28445\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32785\,
            in1 => \N__30761\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31286\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28837\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25744\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32786\,
            in1 => \N__27330\,
            in2 => \_gnd_net_\,
            in3 => \N__28284\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32787\,
            in1 => \N__32376\,
            in2 => \_gnd_net_\,
            in3 => \N__32411\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32030\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28768\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35242\,
            in1 => \N__35606\,
            in2 => \N__31527\,
            in3 => \N__31550\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35609\,
            in1 => \N__35241\,
            in2 => \N__28740\,
            in3 => \N__28769\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__35243\,
            in1 => \N__35607\,
            in2 => \N__28455\,
            in3 => \N__25759\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31519\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__35239\,
            in1 => \N__35608\,
            in2 => \N__31268\,
            in3 => \N__31301\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35605\,
            in1 => \N__35240\,
            in2 => \N__27407\,
            in3 => \N__28511\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28669\,
            in1 => \N__28646\,
            in2 => \_gnd_net_\,
            in3 => \N__30420\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26559\,
            in1 => \N__26537\,
            in2 => \_gnd_net_\,
            in3 => \N__30419\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__25873\,
            in1 => \N__28605\,
            in2 => \N__28584\,
            in3 => \N__28554\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49968\,
            ce => 'H',
            sr => \N__49404\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37126\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49968\,
            ce => 'H',
            sr => \N__49404\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__28604\,
            in1 => \N__25861\,
            in2 => \N__25848\,
            in3 => \N__29149\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49968\,
            ce => 'H',
            sr => \N__49404\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27151\,
            in1 => \N__28945\,
            in2 => \N__26389\,
            in3 => \N__28898\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26284\,
            in1 => \N__26459\,
            in2 => \N__25822\,
            in3 => \N__25807\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29384\,
            in2 => \_gnd_net_\,
            in3 => \N__29351\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30493\,
            in1 => \N__28920\,
            in2 => \_gnd_net_\,
            in3 => \N__28946\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28947\,
            in1 => \_gnd_net_\,
            in2 => \N__25801\,
            in3 => \N__30497\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__29247\,
            sr => \N__49409\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26387\,
            in1 => \_gnd_net_\,
            in2 => \N__30548\,
            in3 => \N__26349\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__29247\,
            sr => \N__49409\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30557\,
            in1 => \N__27121\,
            in2 => \_gnd_net_\,
            in3 => \N__27152\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => \N__29247\,
            sr => \N__49409\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__25954\,
            in1 => \N__25932\,
            in2 => \N__25906\,
            in3 => \N__25891\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__25890\,
            in1 => \N__25953\,
            in2 => \N__25936\,
            in3 => \N__25902\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26489\,
            in1 => \N__26502\,
            in2 => \_gnd_net_\,
            in3 => \N__30437\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30440\,
            in1 => \_gnd_net_\,
            in2 => \N__25909\,
            in3 => \N__26490\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__29252\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29462\,
            in1 => \N__29430\,
            in2 => \_gnd_net_\,
            in3 => \N__30438\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30439\,
            in1 => \_gnd_net_\,
            in2 => \N__25894\,
            in3 => \N__29463\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__29252\,
            sr => \N__49416\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29507\,
            in1 => \N__29539\,
            in2 => \_gnd_net_\,
            in3 => \N__30441\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__29252\,
            sr => \N__49416\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__26233\,
            in1 => \N__26211\,
            in2 => \N__26101\,
            in3 => \N__26086\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26085\,
            in1 => \N__26232\,
            in2 => \N__26215\,
            in3 => \N__26097\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30550\,
            in1 => \N__29360\,
            in2 => \_gnd_net_\,
            in3 => \N__29331\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29361\,
            in1 => \_gnd_net_\,
            in2 => \N__26188\,
            in3 => \N__30553\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__29248\,
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30552\,
            in1 => \N__26173\,
            in2 => \_gnd_net_\,
            in3 => \N__26142\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__29248\,
            sr => \N__49424\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30617\,
            in1 => \N__30573\,
            in2 => \_gnd_net_\,
            in3 => \N__30549\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30551\,
            in1 => \_gnd_net_\,
            in2 => \N__26089\,
            in3 => \N__30618\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__29248\,
            sr => \N__49424\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26077\,
            in1 => \_gnd_net_\,
            in2 => \N__30558\,
            in3 => \N__26038\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26008\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__30534\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30529\,
            in1 => \N__26563\,
            in2 => \_gnd_net_\,
            in3 => \N__26539\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26506\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \N__30535\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30530\,
            in1 => \N__26461\,
            in2 => \_gnd_net_\,
            in3 => \N__26416\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26388\,
            in1 => \N__26350\,
            in2 => \_gnd_net_\,
            in3 => \N__30537\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30528\,
            in1 => \N__26326\,
            in2 => \_gnd_net_\,
            in3 => \N__26302\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26287\,
            in1 => \N__26257\,
            in2 => \_gnd_net_\,
            in3 => \N__30536\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => \N__30103\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__33663\,
            in1 => \N__33636\,
            in2 => \N__26809\,
            in3 => \N__26875\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__26874\,
            in1 => \N__33664\,
            in2 => \N__33640\,
            in3 => \N__26805\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26941\,
            in1 => \N__26913\,
            in2 => \_gnd_net_\,
            in3 => \N__30324\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => \N__30101\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30323\,
            in1 => \N__26866\,
            in2 => \_gnd_net_\,
            in3 => \N__26830\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => \N__30101\,
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__33586\,
            in1 => \N__33609\,
            in2 => \N__26668\,
            in3 => \N__26743\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26742\,
            in1 => \N__33585\,
            in2 => \N__33613\,
            in3 => \N__26664\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30325\,
            in1 => \N__26797\,
            in2 => \_gnd_net_\,
            in3 => \N__26764\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__30100\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26734\,
            in1 => \N__26706\,
            in2 => \_gnd_net_\,
            in3 => \N__30327\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__30100\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30326\,
            in1 => \N__26656\,
            in2 => \_gnd_net_\,
            in3 => \N__26629\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__30100\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__33853\,
            in1 => \N__33873\,
            in2 => \N__27169\,
            in3 => \N__27241\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27240\,
            in1 => \N__33852\,
            in2 => \N__33877\,
            in3 => \N__27165\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27286\,
            in1 => \N__27256\,
            in2 => \_gnd_net_\,
            in3 => \N__30322\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49910\,
            ce => \N__30098\,
            sr => \N__49459\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30321\,
            in1 => \N__27232\,
            in2 => \_gnd_net_\,
            in3 => \N__27207\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49910\,
            ce => \N__30098\,
            sr => \N__49459\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27117\,
            in1 => \N__27153\,
            in2 => \_gnd_net_\,
            in3 => \N__30320\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__33805\,
            in1 => \N__33828\,
            in2 => \N__27019\,
            in3 => \N__27097\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__27096\,
            in1 => \N__33804\,
            in2 => \N__33832\,
            in3 => \N__27015\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27085\,
            in1 => \N__27058\,
            in2 => \_gnd_net_\,
            in3 => \N__30562\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => \N__30096\,
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30561\,
            in1 => \N__27006\,
            in2 => \_gnd_net_\,
            in3 => \N__26971\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => \N__30096\,
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__30021\,
            in1 => \N__30006\,
            in2 => \N__34102\,
            in3 => \N__34129\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31162\,
            in1 => \N__35542\,
            in2 => \N__35147\,
            in3 => \N__31120\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35539\,
            in1 => \N__35013\,
            in2 => \N__31873\,
            in3 => \N__31894\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32775\,
            in1 => \N__27478\,
            in2 => \_gnd_net_\,
            in3 => \N__28241\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35540\,
            in1 => \N__35014\,
            in2 => \N__31729\,
            in3 => \N__31683\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32776\,
            in1 => \N__31778\,
            in2 => \_gnd_net_\,
            in3 => \N__31818\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35544\,
            in1 => \N__35016\,
            in2 => \N__27415\,
            in3 => \N__28522\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31084\,
            in1 => \N__35541\,
            in2 => \N__35146\,
            in3 => \N__30912\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35543\,
            in1 => \N__35015\,
            in2 => \N__32395\,
            in3 => \N__32424\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__28300\,
            in1 => \N__35453\,
            in2 => \N__35072\,
            in3 => \N__27340\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35450\,
            in1 => \N__34901\,
            in2 => \N__30865\,
            in3 => \N__30814\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34895\,
            in1 => \N__35452\,
            in2 => \N__31603\,
            in3 => \N__31641\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35451\,
            in1 => \N__34902\,
            in2 => \N__31369\,
            in3 => \N__31400\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__34896\,
            in1 => \N__35454\,
            in2 => \N__35290\,
            in3 => \N__34645\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35455\,
            in1 => \N__34900\,
            in2 => \N__32074\,
            in3 => \N__32037\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__34893\,
            in1 => \N__35456\,
            in2 => \N__28819\,
            in3 => \N__28864\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35449\,
            in1 => \N__34894\,
            in2 => \N__32155\,
            in3 => \N__32112\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27525\,
            in2 => \N__27508\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32834\,
            in2 => \N__32803\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34921\,
            in2 => \N__31417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30937\,
            in2 => \N__35108\,
            in3 => \N__27706\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34925\,
            in2 => \N__31174\,
            in3 => \N__27691\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27688\,
            in2 => \N__35109\,
            in3 => \N__27670\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34929\,
            in2 => \N__31924\,
            in3 => \N__27655\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31315\,
            in2 => \N__35110\,
            in3 => \N__27637\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34933\,
            in2 => \N__31906\,
            in3 => \N__27619\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32332\,
            in2 => \N__35111\,
            in3 => \N__27598\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34937\,
            in2 => \N__32083\,
            in3 => \N__27586\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32440\,
            in2 => \N__35112\,
            in3 => \N__27853\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34941\,
            in2 => \N__31654\,
            in3 => \N__27835\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27832\,
            in2 => \N__35113\,
            in3 => \N__27814\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34945\,
            in2 => \N__30877\,
            in3 => \N__27799\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31090\,
            in2 => \N__35114\,
            in3 => \N__27781\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35115\,
            in2 => \N__30781\,
            in3 => \N__27763\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31321\,
            in2 => \N__35222\,
            in3 => \N__27742\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35119\,
            in2 => \N__30709\,
            in3 => \N__27724\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31570\,
            in2 => \N__35223\,
            in3 => \N__28015\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35123\,
            in2 => \N__28012\,
            in3 => \N__27991\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32353\,
            in2 => \N__35224\,
            in3 => \N__27976\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35127\,
            in2 => \N__27973\,
            in3 => \N__27946\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34609\,
            in2 => \N__35225\,
            in3 => \N__27931\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35131\,
            in2 => \N__31999\,
            in3 => \N__27916\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35140\,
            in2 => \N__31495\,
            in3 => \N__27901\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35132\,
            in2 => \N__27898\,
            in3 => \N__27871\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35141\,
            in2 => \N__28789\,
            in3 => \N__28126\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35133\,
            in2 => \N__31237\,
            in3 => \N__28111\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35142\,
            in2 => \N__28714\,
            in3 => \N__28093\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35134\,
            in2 => \N__32512\,
            in3 => \N__28075\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__35135\,
            in1 => \N__35601\,
            in2 => \_gnd_net_\,
            in3 => \N__28072\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32851\,
            in2 => \N__32247\,
            in3 => \N__32237\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28057\,
            in2 => \_gnd_net_\,
            in3 => \N__28051\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28048\,
            in2 => \_gnd_net_\,
            in3 => \N__28042\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28039\,
            in2 => \_gnd_net_\,
            in3 => \N__28033\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28261\,
            in2 => \_gnd_net_\,
            in3 => \N__28219\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28216\,
            in2 => \_gnd_net_\,
            in3 => \N__28210\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28207\,
            in2 => \_gnd_net_\,
            in3 => \N__28198\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28195\,
            in2 => \_gnd_net_\,
            in3 => \N__28186\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28183\,
            in2 => \_gnd_net_\,
            in3 => \N__28174\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28171\,
            in2 => \_gnd_net_\,
            in3 => \N__28165\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28162\,
            in2 => \_gnd_net_\,
            in3 => \N__28150\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28147\,
            in2 => \_gnd_net_\,
            in3 => \N__28141\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28393\,
            in2 => \_gnd_net_\,
            in3 => \N__28360\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31042\,
            in2 => \_gnd_net_\,
            in3 => \N__28357\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28354\,
            in2 => \_gnd_net_\,
            in3 => \N__28348\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28345\,
            in2 => \_gnd_net_\,
            in3 => \N__28339\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28336\,
            in2 => \_gnd_net_\,
            in3 => \N__28327\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28324\,
            in2 => \_gnd_net_\,
            in3 => \N__28318\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28315\,
            in2 => \_gnd_net_\,
            in3 => \N__28309\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28306\,
            in2 => \_gnd_net_\,
            in3 => \N__28273\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28270\,
            in2 => \_gnd_net_\,
            in3 => \N__28264\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28528\,
            in2 => \_gnd_net_\,
            in3 => \N__28495\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28492\,
            in2 => \_gnd_net_\,
            in3 => \N__28486\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28483\,
            in2 => \_gnd_net_\,
            in3 => \N__28477\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28474\,
            in2 => \_gnd_net_\,
            in3 => \N__28468\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28465\,
            in2 => \_gnd_net_\,
            in3 => \N__28429\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28426\,
            in2 => \_gnd_net_\,
            in3 => \N__28414\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28411\,
            in2 => \_gnd_net_\,
            in3 => \N__28405\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28402\,
            in2 => \_gnd_net_\,
            in3 => \N__28396\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28867\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__35244\,
            in2 => \N__28863\,
            in3 => \N__28808\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35245\,
            in1 => \N__35611\,
            in2 => \N__28777\,
            in3 => \N__28733\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42013\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49867\,
            ce => 'H',
            sr => \N__49523\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28687\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28667\,
            in1 => \N__28651\,
            in2 => \_gnd_net_\,
            in3 => \N__30424\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49967\,
            ce => \N__30106\,
            sr => \N__49392\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__39996\,
            in1 => \N__28609\,
            in2 => \N__28585\,
            in3 => \N__28555\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49958\,
            ce => 'H',
            sr => \N__49398\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__43448\,
            in1 => \N__43415\,
            in2 => \N__48392\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43799\,
            in1 => \N__43779\,
            in2 => \_gnd_net_\,
            in3 => \N__48362\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__44000\,
            in1 => \N__44024\,
            in2 => \N__48391\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29537\,
            in1 => \N__29517\,
            in2 => \_gnd_net_\,
            in3 => \N__30498\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28907\,
            in1 => \N__28878\,
            in2 => \_gnd_net_\,
            in3 => \N__30490\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30491\,
            in1 => \_gnd_net_\,
            in2 => \N__29302\,
            in3 => \N__28908\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49941\,
            ce => \N__29253\,
            sr => \N__49410\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29395\,
            in1 => \N__29410\,
            in2 => \_gnd_net_\,
            in3 => \N__30492\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49941\,
            ce => \N__29253\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48358\,
            in1 => \N__44159\,
            in2 => \_gnd_net_\,
            in3 => \N__44135\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48570\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28951\,
            in1 => \N__28924\,
            in2 => \_gnd_net_\,
            in3 => \N__30555\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => \N__30105\,
            sr => \N__49417\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28909\,
            in1 => \N__28879\,
            in2 => \_gnd_net_\,
            in3 => \N__30556\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => \N__30105\,
            sr => \N__49417\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30554\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \N__29518\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => \N__30105\,
            sr => \N__49417\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__33561\,
            in1 => \N__29419\,
            in2 => \N__29476\,
            in3 => \N__33903\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__29418\,
            in1 => \N__33562\,
            in2 => \N__33904\,
            in3 => \N__29475\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29464\,
            in1 => \N__29434\,
            in2 => \_gnd_net_\,
            in3 => \N__30435\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => \N__30104\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29393\,
            in1 => \N__29406\,
            in2 => \_gnd_net_\,
            in3 => \N__30433\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__30434\,
            in1 => \N__29394\,
            in2 => \N__29365\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => \N__30104\,
            sr => \N__49425\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29362\,
            in1 => \N__29332\,
            in2 => \_gnd_net_\,
            in3 => \N__30436\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => \N__30104\,
            sr => \N__49425\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29308\,
            in2 => \N__29320\,
            in3 => \N__41538\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29674\,
            in2 => \N__29668\,
            in3 => \N__33378\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29659\,
            in2 => \N__29647\,
            in3 => \N__33360\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29638\,
            in2 => \N__29629\,
            in3 => \N__33540\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29620\,
            in2 => \N__29614\,
            in3 => \N__33526\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29593\,
            in2 => \N__29602\,
            in3 => \N__33507\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29578\,
            in2 => \N__29587\,
            in3 => \N__33492\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29563\,
            in2 => \N__29572\,
            in3 => \N__33477\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29557\,
            in2 => \N__29548\,
            in3 => \N__33463\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33445\,
            in1 => \N__29809\,
            in2 => \N__29821\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29791\,
            in2 => \N__29803\,
            in3 => \N__33426\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29785\,
            in2 => \N__29776\,
            in3 => \N__33411\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \N__29752\,
            in3 => \N__33708\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29743\,
            in2 => \N__29734\,
            in3 => \N__33693\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29725\,
            in2 => \N__29716\,
            in3 => \N__33678\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29707\,
            in2 => \N__29701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29692\,
            in2 => \N__29686\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29896\,
            in2 => \N__29887\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29875\,
            in2 => \N__29866\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29854\,
            in2 => \N__29848\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30682\,
            in2 => \N__29830\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30067\,
            in2 => \N__30034\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29839\,
            in2 => \N__29992\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29833\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__33783\,
            in1 => \N__30696\,
            in2 => \N__33766\,
            in3 => \N__30628\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__30627\,
            in1 => \N__33761\,
            in2 => \N__30700\,
            in3 => \N__33782\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30676\,
            in1 => \N__30646\,
            in2 => \_gnd_net_\,
            in3 => \N__30559\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => \N__30099\,
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30619\,
            in1 => \N__30580\,
            in2 => \_gnd_net_\,
            in3 => \N__30560\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => \N__30099\,
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__30042\,
            in1 => \N__33722\,
            in2 => \N__30061\,
            in3 => \N__33743\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__33723\,
            in1 => \N__30057\,
            in2 => \N__33745\,
            in3 => \N__30043\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__30025\,
            in1 => \N__34097\,
            in2 => \N__30007\,
            in3 => \N__34127\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29979\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49472\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29953\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49472\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29925\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49472\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31030\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49472\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35186\,
            in1 => \N__35423\,
            in2 => \N__30987\,
            in3 => \N__30957\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32188\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__32878\,
            sr => \N__49479\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35187\,
            in1 => \N__35424\,
            in2 => \N__30988\,
            in3 => \N__30958\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35422\,
            in1 => \N__35188\,
            in2 => \N__31482\,
            in3 => \N__31441\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35426\,
            in1 => \N__35227\,
            in2 => \N__30913\,
            in3 => \N__31080\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35228\,
            in1 => \N__35427\,
            in2 => \N__30864\,
            in3 => \N__30813\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35429\,
            in1 => \N__35226\,
            in2 => \N__30772\,
            in3 => \N__30733\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35430\,
            in1 => \N__35229\,
            in2 => \N__31564\,
            in3 => \N__31528\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35425\,
            in1 => \N__35231\,
            in2 => \N__31483\,
            in3 => \N__31437\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__35230\,
            in1 => \N__35428\,
            in2 => \N__31405\,
            in3 => \N__31365\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35497\,
            in1 => \N__35175\,
            in2 => \N__31782\,
            in3 => \N__31819\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31306\,
            in1 => \N__35501\,
            in2 => \N__35234\,
            in3 => \N__31270\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31228\,
            in1 => \N__35496\,
            in2 => \N__35233\,
            in3 => \N__31201\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35499\,
            in1 => \N__35176\,
            in2 => \N__31161\,
            in3 => \N__31119\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31072\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35498\,
            in1 => \N__35171\,
            in2 => \N__32151\,
            in3 => \N__32111\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__35177\,
            in1 => \N__32067\,
            in2 => \N__32041\,
            in3 => \N__35500\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__35562\,
            in1 => \N__35215\,
            in2 => \N__31990\,
            in3 => \N__31960\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35218\,
            in1 => \N__35564\,
            in2 => \N__31872\,
            in3 => \N__31887\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__31886\,
            in1 => \N__32704\,
            in2 => \_gnd_net_\,
            in3 => \N__31865\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__35216\,
            in1 => \N__35563\,
            in2 => \N__31814\,
            in3 => \N__31786\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__35566\,
            in1 => \N__35219\,
            in2 => \N__31722\,
            in3 => \N__31682\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__35221\,
            in1 => \N__35567\,
            in2 => \N__31642\,
            in3 => \N__31598\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__35565\,
            in1 => \N__32494\,
            in2 => \N__32470\,
            in3 => \N__35217\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__35220\,
            in1 => \N__35568\,
            in2 => \N__32428\,
            in3 => \N__32391\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__32274\,
            in1 => \N__35569\,
            in2 => \N__32305\,
            in3 => \N__35164\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35570\,
            in1 => \N__32304\,
            in2 => \N__35232\,
            in3 => \N__32275\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35571\,
            in2 => \_gnd_net_\,
            in3 => \N__35163\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32300\,
            in1 => \N__32683\,
            in2 => \_gnd_net_\,
            in3 => \N__32273\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32939\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__32940\,
            in1 => \_gnd_net_\,
            in2 => \N__32218\,
            in3 => \N__32682\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32184\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__32875\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32977\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__32875\,
            sr => \N__49498\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__35536\,
            in1 => \N__32643\,
            in2 => \N__32839\,
            in3 => \N__32631\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32905\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49873\,
            ce => \N__32874\,
            sr => \N__49502\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32629\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__32632\,
            in1 => \N__35537\,
            in2 => \N__32647\,
            in3 => \N__32838\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__32684\,
            in1 => \N__32642\,
            in2 => \_gnd_net_\,
            in3 => \N__32630\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__35538\,
            in1 => \N__35236\,
            in2 => \N__32599\,
            in3 => \N__32534\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34527\,
            in2 => \_gnd_net_\,
            in3 => \N__34593\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__34468\,
            in1 => \N__34495\,
            in2 => \N__32497\,
            in3 => \N__34564\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35706\,
            in1 => \N__35733\,
            in2 => \_gnd_net_\,
            in3 => \N__35759\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__35787\,
            in1 => \N__33007\,
            in2 => \N__33001\,
            in3 => \N__34437\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33071\,
            in1 => \N__34592\,
            in2 => \_gnd_net_\,
            in3 => \N__32998\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_26_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_1_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33067\,
            in1 => \N__34556\,
            in2 => \_gnd_net_\,
            in3 => \N__32995\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_2_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33072\,
            in1 => \N__34526\,
            in2 => \_gnd_net_\,
            in3 => \N__32992\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_3_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33068\,
            in1 => \N__34493\,
            in2 => \_gnd_net_\,
            in3 => \N__32989\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_4_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33073\,
            in1 => \N__34466\,
            in2 => \_gnd_net_\,
            in3 => \N__32986\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_5_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33069\,
            in1 => \N__34436\,
            in2 => \_gnd_net_\,
            in3 => \N__32983\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_6_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33074\,
            in1 => \N__35786\,
            in2 => \_gnd_net_\,
            in3 => \N__32980\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_7_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33070\,
            in1 => \N__35760\,
            in2 => \_gnd_net_\,
            in3 => \N__33082\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49517\
        );

    \pwm_generator_inst.counter_8_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33076\,
            in1 => \N__35732\,
            in2 => \_gnd_net_\,
            in3 => \N__33079\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__49865\,
            ce => 'H',
            sr => \N__49521\
        );

    \pwm_generator_inst.counter_9_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35705\,
            in1 => \N__33075\,
            in2 => \_gnd_net_\,
            in3 => \N__33034\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49865\,
            ce => 'H',
            sr => \N__49521\
        );

    \GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_red_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36009\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49978\,
            ce => \N__36462\,
            sr => \N__49385\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35988\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49978\,
            ce => \N__36462\,
            sr => \N__49385\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33320\,
            in1 => \N__36005\,
            in2 => \_gnd_net_\,
            in3 => \N__33016\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33315\,
            in1 => \N__35984\,
            in2 => \_gnd_net_\,
            in3 => \N__33013\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33321\,
            in1 => \N__35961\,
            in2 => \_gnd_net_\,
            in3 => \N__33010\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33316\,
            in1 => \N__35937\,
            in2 => \_gnd_net_\,
            in3 => \N__33109\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33322\,
            in1 => \N__35913\,
            in2 => \_gnd_net_\,
            in3 => \N__33106\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33317\,
            in1 => \N__35889\,
            in2 => \_gnd_net_\,
            in3 => \N__33103\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33319\,
            in1 => \N__35865\,
            in2 => \_gnd_net_\,
            in3 => \N__33100\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33318\,
            in1 => \N__35841\,
            in2 => \_gnd_net_\,
            in3 => \N__33097\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49969\,
            ce => \N__33187\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33311\,
            in1 => \N__36198\,
            in2 => \_gnd_net_\,
            in3 => \N__33094\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33296\,
            in1 => \N__36174\,
            in2 => \_gnd_net_\,
            in3 => \N__33091\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33308\,
            in1 => \N__36150\,
            in2 => \_gnd_net_\,
            in3 => \N__33088\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__36126\,
            in2 => \_gnd_net_\,
            in3 => \N__33085\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33309\,
            in1 => \N__36102\,
            in2 => \_gnd_net_\,
            in3 => \N__33136\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33294\,
            in1 => \N__36078\,
            in2 => \_gnd_net_\,
            in3 => \N__33133\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33310\,
            in1 => \N__36054\,
            in2 => \_gnd_net_\,
            in3 => \N__33130\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33295\,
            in1 => \N__36030\,
            in2 => \_gnd_net_\,
            in3 => \N__33127\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49960\,
            ce => \N__33182\,
            sr => \N__49399\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33297\,
            in1 => \N__36387\,
            in2 => \_gnd_net_\,
            in3 => \N__33124\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33301\,
            in1 => \N__36363\,
            in2 => \_gnd_net_\,
            in3 => \N__33121\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33298\,
            in1 => \N__36343\,
            in2 => \_gnd_net_\,
            in3 => \N__33118\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33302\,
            in1 => \N__36321\,
            in2 => \_gnd_net_\,
            in3 => \N__33115\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33299\,
            in1 => \N__36299\,
            in2 => \_gnd_net_\,
            in3 => \N__33112\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33303\,
            in1 => \N__36273\,
            in2 => \_gnd_net_\,
            in3 => \N__33346\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33300\,
            in1 => \N__36249\,
            in2 => \_gnd_net_\,
            in3 => \N__33343\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33304\,
            in1 => \N__36225\,
            in2 => \_gnd_net_\,
            in3 => \N__33340\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49951\,
            ce => \N__33181\,
            sr => \N__49405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33312\,
            in1 => \N__36582\,
            in2 => \_gnd_net_\,
            in3 => \N__33337\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33305\,
            in1 => \N__36558\,
            in2 => \_gnd_net_\,
            in3 => \N__33334\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__36522\,
            in2 => \_gnd_net_\,
            in3 => \N__33331\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33306\,
            in1 => \N__36486\,
            in2 => \_gnd_net_\,
            in3 => \N__33328\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33314\,
            in1 => \N__36538\,
            in2 => \_gnd_net_\,
            in3 => \N__33325\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33307\,
            in1 => \N__36502\,
            in2 => \_gnd_net_\,
            in3 => \N__33190\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => \N__33186\,
            sr => \N__49411\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__33397\,
            in1 => \N__39829\,
            in2 => \N__39805\,
            in3 => \N__33388\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41518\,
            in1 => \N__41489\,
            in2 => \_gnd_net_\,
            in3 => \N__48398\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => \N__45840\,
            sr => \N__49418\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48397\,
            in1 => \N__41431\,
            in2 => \_gnd_net_\,
            in3 => \N__41407\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => \N__45840\,
            sr => \N__49418\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__33396\,
            in1 => \N__39828\,
            in2 => \N__39804\,
            in3 => \N__33387\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47524\,
            in1 => \N__47500\,
            in2 => \_gnd_net_\,
            in3 => \N__48399\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => \N__45840\,
            sr => \N__49418\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__36645\,
            in1 => \N__39687\,
            in2 => \N__39724\,
            in3 => \N__36633\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41539\,
            in2 => \N__36622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41230\,
            in1 => \N__33379\,
            in2 => \_gnd_net_\,
            in3 => \N__33367\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__41260\,
            in1 => \N__36607\,
            in2 => \N__33364\,
            in3 => \N__33349\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41231\,
            in1 => \N__33541\,
            in2 => \_gnd_net_\,
            in3 => \N__33529\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41261\,
            in1 => \N__33525\,
            in2 => \_gnd_net_\,
            in3 => \N__33511\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41232\,
            in1 => \N__33508\,
            in2 => \_gnd_net_\,
            in3 => \N__33496\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41262\,
            in1 => \N__33493\,
            in2 => \_gnd_net_\,
            in3 => \N__33481\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41233\,
            in1 => \N__33478\,
            in2 => \_gnd_net_\,
            in3 => \N__33466\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41255\,
            in1 => \N__33462\,
            in2 => \_gnd_net_\,
            in3 => \N__33448\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41256\,
            in1 => \N__33444\,
            in2 => \_gnd_net_\,
            in3 => \N__33430\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41252\,
            in1 => \N__33427\,
            in2 => \_gnd_net_\,
            in3 => \N__33415\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41257\,
            in1 => \N__33412\,
            in2 => \_gnd_net_\,
            in3 => \N__33400\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41253\,
            in1 => \N__33709\,
            in2 => \_gnd_net_\,
            in3 => \N__33697\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41258\,
            in1 => \N__33694\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41254\,
            in1 => \N__33679\,
            in2 => \_gnd_net_\,
            in3 => \N__33667\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41259\,
            in1 => \N__33657\,
            in2 => \_gnd_net_\,
            in3 => \N__33643\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49915\,
            ce => 'H',
            sr => \N__49433\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41240\,
            in1 => \N__33630\,
            in2 => \_gnd_net_\,
            in3 => \N__33616\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41244\,
            in1 => \N__33603\,
            in2 => \_gnd_net_\,
            in3 => \N__33589\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41241\,
            in1 => \N__33579\,
            in2 => \_gnd_net_\,
            in3 => \N__33565\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41245\,
            in1 => \N__33560\,
            in2 => \_gnd_net_\,
            in3 => \N__33544\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41242\,
            in1 => \N__33894\,
            in2 => \_gnd_net_\,
            in3 => \N__33880\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41246\,
            in1 => \N__33872\,
            in2 => \_gnd_net_\,
            in3 => \N__33856\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41243\,
            in1 => \N__33851\,
            in2 => \_gnd_net_\,
            in3 => \N__33835\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41247\,
            in1 => \N__33822\,
            in2 => \_gnd_net_\,
            in3 => \N__33808\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49911\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41248\,
            in1 => \N__33803\,
            in2 => \_gnd_net_\,
            in3 => \N__33787\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41237\,
            in1 => \N__33784\,
            in2 => \_gnd_net_\,
            in3 => \N__33769\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41249\,
            in1 => \N__33765\,
            in2 => \_gnd_net_\,
            in3 => \N__33748\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41238\,
            in1 => \N__33744\,
            in2 => \_gnd_net_\,
            in3 => \N__33727\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41250\,
            in1 => \N__33724\,
            in2 => \_gnd_net_\,
            in3 => \N__34132\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41239\,
            in1 => \N__34128\,
            in2 => \_gnd_net_\,
            in3 => \N__34108\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41251\,
            in1 => \N__34098\,
            in2 => \_gnd_net_\,
            in3 => \N__34105\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49905\,
            ce => 'H',
            sr => \N__49451\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34078\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34048\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33994\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33964\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49896\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33936\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49896\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34411\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49896\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34384\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49896\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34353\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49473\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34329\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49473\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34300\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49473\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34272\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49885\,
            ce => 'H',
            sr => \N__49480\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34242\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49885\,
            ce => 'H',
            sr => \N__49480\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34209\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49885\,
            ce => 'H',
            sr => \N__49480\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34176\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49885\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst1.S2_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49880\,
            ce => 'H',
            sr => \N__49485\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35643\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49880\,
            ce => 'H',
            sr => \N__49485\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__35572\,
            in1 => \N__35279\,
            in2 => \N__35235\,
            in3 => \N__34638\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34570\,
            in2 => \N__38857\,
            in3 => \N__34597\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38557\,
            in2 => \N__34540\,
            in3 => \N__34563\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38887\,
            in2 => \N__34504\,
            in3 => \N__34531\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34474\,
            in2 => \N__38572\,
            in3 => \N__34494\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34467\,
            in1 => \N__38587\,
            in2 => \N__34447\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34438\,
            in1 => \N__34417\,
            in2 => \N__38542\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35788\,
            in1 => \N__35767\,
            in2 => \N__38602\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35761\,
            in1 => \N__35740\,
            in2 => \N__38872\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35713\,
            in2 => \N__38839\,
            in3 => \N__35734\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35683\,
            in2 => \N__35800\,
            in3 => \N__35707\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35677\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49508\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38830\,
            in2 => \N__44989\,
            in3 => \N__44976\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44866\,
            in2 => \_gnd_net_\,
            in3 => \N__35650\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38818\,
            in2 => \_gnd_net_\,
            in3 => \N__35647\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38824\,
            in2 => \_gnd_net_\,
            in3 => \N__35824\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38812\,
            in2 => \_gnd_net_\,
            in3 => \N__35821\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42169\,
            in2 => \_gnd_net_\,
            in3 => \N__35818\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43219\,
            in2 => \_gnd_net_\,
            in3 => \N__35815\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38926\,
            in2 => \_gnd_net_\,
            in3 => \N__35812\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43231\,
            in2 => \_gnd_net_\,
            in3 => \N__35809\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_13_27_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__45166\,
            in1 => \N__40396\,
            in2 => \N__44992\,
            in3 => \N__35806\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__49051\,
            in1 => \N__47848\,
            in2 => \N__35803\,
            in3 => \N__42312\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44091\,
            in1 => \N__44069\,
            in2 => \_gnd_net_\,
            in3 => \N__48329\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45536\,
            in1 => \N__45509\,
            in2 => \_gnd_net_\,
            in3 => \N__48348\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35960\,
            in2 => \N__36010\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35936\,
            in2 => \N__35989\,
            in3 => \N__35968\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35912\,
            in2 => \N__35965\,
            in3 => \N__35944\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35888\,
            in2 => \N__35941\,
            in3 => \N__35920\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35864\,
            in2 => \N__35917\,
            in3 => \N__35896\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35840\,
            in2 => \N__35893\,
            in3 => \N__35872\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36197\,
            in2 => \N__35869\,
            in3 => \N__35848\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36173\,
            in2 => \N__35845\,
            in3 => \N__36205\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49979\,
            ce => \N__36463\,
            sr => \N__49386\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36149\,
            in2 => \N__36202\,
            in3 => \N__36181\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36125\,
            in2 => \N__36178\,
            in3 => \N__36157\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36101\,
            in2 => \N__36154\,
            in3 => \N__36133\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36077\,
            in2 => \N__36130\,
            in3 => \N__36109\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36053\,
            in2 => \N__36106\,
            in3 => \N__36085\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36029\,
            in2 => \N__36082\,
            in3 => \N__36061\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36386\,
            in2 => \N__36058\,
            in3 => \N__36037\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36362\,
            in2 => \N__36034\,
            in3 => \N__36013\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49970\,
            ce => \N__36461\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36341\,
            in2 => \N__36391\,
            in3 => \N__36370\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36320\,
            in2 => \N__36367\,
            in3 => \N__36346\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36342\,
            in2 => \N__36300\,
            in3 => \N__36328\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36272\,
            in2 => \N__36325\,
            in3 => \N__36304\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36248\,
            in2 => \N__36301\,
            in3 => \N__36280\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36224\,
            in2 => \N__36277\,
            in3 => \N__36256\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36581\,
            in2 => \N__36253\,
            in3 => \N__36232\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36557\,
            in2 => \N__36229\,
            in3 => \N__36208\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49961\,
            ce => \N__36447\,
            sr => \N__49400\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36521\,
            in2 => \N__36586\,
            in3 => \N__36565\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49952\,
            ce => \N__36460\,
            sr => \N__49406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36485\,
            in2 => \N__36562\,
            in3 => \N__36541\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49952\,
            ce => \N__36460\,
            sr => \N__49406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36537\,
            in2 => \N__36526\,
            in3 => \N__36505\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49952\,
            ce => \N__36460\,
            sr => \N__49406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36501\,
            in2 => \N__36490\,
            in3 => \N__36469\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49952\,
            ce => \N__36460\,
            sr => \N__49406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36466\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => \N__36460\,
            sr => \N__49406\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__39748\,
            in1 => \N__39771\,
            in2 => \N__36403\,
            in3 => \N__36655\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__36654\,
            in1 => \N__39747\,
            in2 => \N__39775\,
            in3 => \N__36399\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41879\,
            in1 => \N__48393\,
            in2 => \_gnd_net_\,
            in3 => \N__41898\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48395\,
            in1 => \_gnd_net_\,
            in2 => \N__36406\,
            in3 => \N__41880\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => \N__45844\,
            sr => \N__49412\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48394\,
            in1 => \N__46168\,
            in2 => \_gnd_net_\,
            in3 => \N__46146\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => \N__45844\,
            sr => \N__49412\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48613\,
            in1 => \N__48649\,
            in2 => \_gnd_net_\,
            in3 => \N__48396\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => \N__45844\,
            sr => \N__49412\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__36646\,
            in1 => \N__39723\,
            in2 => \N__39691\,
            in3 => \N__36634\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41582\,
            in2 => \_gnd_net_\,
            in3 => \N__41553\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41303\,
            in2 => \_gnd_net_\,
            in3 => \N__36771\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36610\,
            in3 => \N__41583\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__36793\,
            in1 => \N__39568\,
            in2 => \N__36601\,
            in3 => \N__39585\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47632\,
            in1 => \N__47593\,
            in2 => \_gnd_net_\,
            in3 => \N__48383\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => \N__45835\,
            sr => \N__49427\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__36792\,
            in1 => \N__39567\,
            in2 => \N__36600\,
            in3 => \N__39584\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47722\,
            in1 => \N__47689\,
            in2 => \_gnd_net_\,
            in3 => \N__48382\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => \N__45835\,
            sr => \N__49427\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44035\,
            in1 => \N__44001\,
            in2 => \_gnd_net_\,
            in3 => \N__48384\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => \N__45835\,
            sr => \N__49427\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__41770\,
            in1 => \N__41335\,
            in2 => \N__39407\,
            in3 => \N__45828\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__41295\,
            in1 => \N__36780\,
            in2 => \_gnd_net_\,
            in3 => \N__42147\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000111010"
        )
    port map (
            in0 => \N__36781\,
            in1 => \N__41296\,
            in2 => \N__36784\,
            in3 => \N__36767\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42148\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__36772\,
            in1 => \N__40354\,
            in2 => \N__41307\,
            in3 => \N__41578\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36741\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36715\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36685\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49452\
        );

    \phase_controller_inst1.state_2_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__41717\,
            in1 => \N__42443\,
            in2 => \N__40018\,
            in3 => \N__40035\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49452\
        );

    \phase_controller_inst1.start_timer_hc_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__41730\,
            in1 => \N__44739\,
            in2 => \N__37115\,
            in3 => \N__39658\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49452\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46695\,
            in2 => \N__39946\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37093\,
            in2 => \N__37084\,
            in3 => \N__37045\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37042\,
            in2 => \N__37036\,
            in3 => \N__36985\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36982\,
            in2 => \N__36976\,
            in3 => \N__36925\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39952\,
            in2 => \N__36922\,
            in3 => \N__36865\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36862\,
            in2 => \N__36853\,
            in3 => \N__36796\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37615\,
            in2 => \N__37606\,
            in3 => \N__37555\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37552\,
            in2 => \N__37546\,
            in3 => \N__37498\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37495\,
            in2 => \N__37489\,
            in3 => \N__37438\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37435\,
            in2 => \N__37378\,
            in3 => \N__37366\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37363\,
            in2 => \N__37351\,
            in3 => \N__37306\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37303\,
            in2 => \N__37294\,
            in3 => \N__37243\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37240\,
            in2 => \N__37234\,
            in3 => \N__37183\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37180\,
            in2 => \N__37174\,
            in3 => \N__37129\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38062\,
            in2 => \N__38047\,
            in3 => \N__37999\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37996\,
            in2 => \N__37990\,
            in3 => \N__37942\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37939\,
            in2 => \N__37933\,
            in3 => \N__37891\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37888\,
            in2 => \N__37849\,
            in3 => \N__37840\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37837\,
            in2 => \N__37795\,
            in3 => \N__37783\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37780\,
            in2 => \N__37774\,
            in3 => \N__37723\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37720\,
            in2 => \N__37711\,
            in3 => \N__37675\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37672\,
            in2 => \N__37666\,
            in3 => \N__37618\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38533\,
            in2 => \N__38521\,
            in3 => \N__38473\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38470\,
            in2 => \N__38461\,
            in3 => \N__38410\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38407\,
            in2 => \N__38398\,
            in3 => \N__38359\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38356\,
            in2 => \N__38347\,
            in3 => \N__38299\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38296\,
            in2 => \N__38281\,
            in3 => \N__38233\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38230\,
            in2 => \N__38191\,
            in3 => \N__38182\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38179\,
            in2 => \N__38173\,
            in3 => \N__38128\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38125\,
            in2 => \N__38110\,
            in3 => \N__38806\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38617\,
            in1 => \N__38801\,
            in2 => \_gnd_net_\,
            in3 => \N__38635\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38632\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => 'H',
            sr => \N__49481\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40383\,
            in2 => \_gnd_net_\,
            in3 => \N__40355\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__49046\,
            in1 => \N__47843\,
            in2 => \N__38611\,
            in3 => \N__42310\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__47841\,
            in1 => \N__38593\,
            in2 => \N__42359\,
            in3 => \N__49044\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__49043\,
            in1 => \N__47840\,
            in2 => \N__38581\,
            in3 => \N__42305\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__47838\,
            in1 => \N__38563\,
            in2 => \N__42357\,
            in3 => \N__49041\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__49045\,
            in1 => \N__47842\,
            in2 => \N__38551\,
            in3 => \N__42309\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__47839\,
            in1 => \N__38893\,
            in2 => \N__42358\,
            in3 => \N__49042\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__49047\,
            in1 => \N__47844\,
            in2 => \N__38881\,
            in3 => \N__42311\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__47818\,
            in1 => \N__38863\,
            in2 => \N__42356\,
            in3 => \N__49016\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__49017\,
            in1 => \N__47819\,
            in2 => \N__42360\,
            in3 => \N__38845\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__46678\,
            in1 => \N__46654\,
            in2 => \N__44990\,
            in3 => \N__45004\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__44984\,
            in1 => \N__45316\,
            in2 => \N__42913\,
            in3 => \N__45340\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__44983\,
            in1 => \N__44824\,
            in2 => \N__44851\,
            in3 => \N__42193\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__45304\,
            in1 => \N__45280\,
            in2 => \N__44991\,
            in3 => \N__42160\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40800\,
            in2 => \_gnd_net_\,
            in3 => \N__45234\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__40801\,
            in1 => \N__45220\,
            in2 => \N__38929\,
            in3 => \N__44985\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42502\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49868\,
            ce => 'H',
            sr => \N__49518\
        );

    \CONSTANT_ONE_LUT4_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43739\,
            in1 => \N__43723\,
            in2 => \_gnd_net_\,
            in3 => \N__48331\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50010\,
            ce => \N__45824\,
            sr => \N__49376\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48330\,
            in1 => \N__44087\,
            in2 => \_gnd_net_\,
            in3 => \N__44070\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50010\,
            ce => \N__45824\,
            sr => \N__49376\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43564\,
            in1 => \N__43187\,
            in2 => \_gnd_net_\,
            in3 => \N__48350\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__45827\,
            sr => \N__49378\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47358\,
            in1 => \N__47387\,
            in2 => \_gnd_net_\,
            in3 => \N__48351\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__45827\,
            sr => \N__49378\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48349\,
            in1 => \N__43205\,
            in2 => \_gnd_net_\,
            in3 => \N__43597\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50003\,
            ce => \N__45827\,
            sr => \N__49378\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__39636\,
            in1 => \N__38901\,
            in2 => \N__39613\,
            in3 => \N__38938\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__38937\,
            in1 => \N__39637\,
            in2 => \N__38905\,
            in3 => \N__39612\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47386\,
            in1 => \N__43660\,
            in2 => \N__47693\,
            in3 => \N__47323\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47594\,
            in1 => \N__41878\,
            in2 => \N__48623\,
            in3 => \N__41485\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45399\,
            in1 => \N__45369\,
            in2 => \_gnd_net_\,
            in3 => \N__48319\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43706\,
            in1 => \N__47224\,
            in2 => \N__47180\,
            in3 => \N__43846\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48324\,
            in1 => \N__43801\,
            in2 => \_gnd_net_\,
            in3 => \N__43771\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45537\,
            in1 => \N__45502\,
            in2 => \_gnd_net_\,
            in3 => \N__48326\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48323\,
            in1 => \N__45901\,
            in2 => \_gnd_net_\,
            in3 => \N__45928\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45397\,
            in1 => \N__45365\,
            in2 => \_gnd_net_\,
            in3 => \N__48327\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48322\,
            in1 => \N__45467\,
            in2 => \_gnd_net_\,
            in3 => \N__45442\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48321\,
            in1 => \N__43690\,
            in2 => \_gnd_net_\,
            in3 => \N__43661\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43825\,
            in1 => \N__43853\,
            in2 => \_gnd_net_\,
            in3 => \N__48325\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49980\,
            ce => \N__45826\,
            sr => \N__49387\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39037\,
            in2 => \N__41104\,
            in3 => \N__39408\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40987\,
            in2 => \N__39031\,
            in3 => \N__39382\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39013\,
            in2 => \N__39022\,
            in3 => \N__39364\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39007\,
            in2 => \N__39001\,
            in3 => \N__39346\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38989\,
            in2 => \N__38983\,
            in3 => \N__39328\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39310\,
            in1 => \N__38971\,
            in2 => \N__38965\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38956\,
            in2 => \N__38947\,
            in3 => \N__39292\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39157\,
            in2 => \N__39145\,
            in3 => \N__39274\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39136\,
            in2 => \N__39127\,
            in3 => \N__39547\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41116\,
            in2 => \N__39118\,
            in3 => \N__39529\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39097\,
            in2 => \N__39109\,
            in3 => \N__39511\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39091\,
            in2 => \N__41095\,
            in3 => \N__39493\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39475\,
            in1 => \N__39073\,
            in2 => \N__39085\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41359\,
            in2 => \N__39067\,
            in3 => \N__39457\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39058\,
            in2 => \N__39049\,
            in3 => \N__39436\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40813\,
            in2 => \N__40876\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40909\,
            in2 => \N__40981\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40996\,
            in2 => \N__41083\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39256\,
            in2 => \N__39247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39232\,
            in2 => \N__39223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39211\,
            in2 => \N__39202\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39190\,
            in2 => \N__39184\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39175\,
            in2 => \N__39169\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39415\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41341\,
            in2 => \N__39412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45773\,
            in1 => \N__39381\,
            in2 => \_gnd_net_\,
            in3 => \N__39367\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__45832\,
            in1 => \N__39363\,
            in2 => \N__41317\,
            in3 => \N__39349\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45774\,
            in1 => \N__39345\,
            in2 => \_gnd_net_\,
            in3 => \N__39331\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45833\,
            in1 => \N__39327\,
            in2 => \_gnd_net_\,
            in3 => \N__39313\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45775\,
            in1 => \N__39309\,
            in2 => \_gnd_net_\,
            in3 => \N__39295\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45834\,
            in1 => \N__39291\,
            in2 => \_gnd_net_\,
            in3 => \N__39277\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45776\,
            in1 => \N__39273\,
            in2 => \_gnd_net_\,
            in3 => \N__39259\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49946\,
            ce => 'H',
            sr => \N__49413\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45780\,
            in1 => \N__39546\,
            in2 => \_gnd_net_\,
            in3 => \N__39532\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45769\,
            in1 => \N__39528\,
            in2 => \_gnd_net_\,
            in3 => \N__39514\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45777\,
            in1 => \N__39510\,
            in2 => \_gnd_net_\,
            in3 => \N__39496\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45770\,
            in1 => \N__39492\,
            in2 => \_gnd_net_\,
            in3 => \N__39478\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45778\,
            in1 => \N__39474\,
            in2 => \_gnd_net_\,
            in3 => \N__39460\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45771\,
            in1 => \N__39453\,
            in2 => \_gnd_net_\,
            in3 => \N__39439\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45779\,
            in1 => \N__39435\,
            in2 => \_gnd_net_\,
            in3 => \N__39421\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45772\,
            in1 => \N__40848\,
            in2 => \_gnd_net_\,
            in3 => \N__39418\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49934\,
            ce => 'H',
            sr => \N__49419\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45757\,
            in1 => \N__40827\,
            in2 => \_gnd_net_\,
            in3 => \N__39652\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45781\,
            in1 => \N__40938\,
            in2 => \_gnd_net_\,
            in3 => \N__39649\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45758\,
            in1 => \N__40962\,
            in2 => \_gnd_net_\,
            in3 => \N__39646\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45782\,
            in1 => \N__41024\,
            in2 => \_gnd_net_\,
            in3 => \N__39643\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45759\,
            in1 => \N__41049\,
            in2 => \_gnd_net_\,
            in3 => \N__39640\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45783\,
            in1 => \N__39630\,
            in2 => \_gnd_net_\,
            in3 => \N__39616\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45760\,
            in1 => \N__39603\,
            in2 => \_gnd_net_\,
            in3 => \N__39589\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45784\,
            in1 => \N__39586\,
            in2 => \_gnd_net_\,
            in3 => \N__39571\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49926\,
            ce => 'H',
            sr => \N__49428\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45753\,
            in1 => \N__39566\,
            in2 => \_gnd_net_\,
            in3 => \N__39550\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45814\,
            in1 => \N__39822\,
            in2 => \_gnd_net_\,
            in3 => \N__39808\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45754\,
            in1 => \N__39792\,
            in2 => \_gnd_net_\,
            in3 => \N__39778\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45815\,
            in1 => \N__39765\,
            in2 => \_gnd_net_\,
            in3 => \N__39751\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45755\,
            in1 => \N__39741\,
            in2 => \_gnd_net_\,
            in3 => \N__39727\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45816\,
            in1 => \N__39713\,
            in2 => \_gnd_net_\,
            in3 => \N__39697\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__45756\,
            in1 => \N__39680\,
            in2 => \_gnd_net_\,
            in3 => \N__39694\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.stoper_tr.running_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001110100"
        )
    port map (
            in0 => \N__41801\,
            in1 => \N__41760\,
            in2 => \N__41818\,
            in3 => \N__41842\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49435\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__40014\,
            in1 => \N__41678\,
            in2 => \N__40036\,
            in3 => \N__41617\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41718\,
            in2 => \_gnd_net_\,
            in3 => \N__42423\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40031\,
            in2 => \_gnd_net_\,
            in3 => \N__40013\,
            lcout => \phase_controller_inst1.state_RNIE87FZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39982\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46696\,
            in2 => \_gnd_net_\,
            in3 => \N__39932\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40047\,
            in1 => \N__40200\,
            in2 => \N__40231\,
            in3 => \N__40071\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39864\,
            in2 => \_gnd_net_\,
            in3 => \N__39883\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40171\,
            in1 => \N__39874\,
            in2 => \N__39886\,
            in3 => \N__40186\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39882\,
            in1 => \N__39853\,
            in2 => \N__39844\,
            in3 => \N__40216\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39873\,
            in1 => \N__39865\,
            in2 => \N__39856\,
            in3 => \N__40117\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39852\,
            in2 => \_gnd_net_\,
            in3 => \N__39840\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40227\,
            in1 => \N__40212\,
            in2 => \N__40201\,
            in3 => \N__40179\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__40180\,
            in1 => \_gnd_net_\,
            in2 => \N__40135\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41967\,
            in1 => \N__40167\,
            in2 => \N__40156\,
            in3 => \N__41913\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40153\,
            in1 => \N__40087\,
            in2 => \N__40147\,
            in3 => \N__40144\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40098\,
            in1 => \N__40131\,
            in2 => \N__40111\,
            in3 => \N__40123\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41931\,
            in2 => \_gnd_net_\,
            in3 => \N__41949\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40107\,
            in1 => \N__40056\,
            in2 => \N__40099\,
            in3 => \N__40080\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40081\,
            in1 => \N__40072\,
            in2 => \N__40060\,
            in3 => \N__40048\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__42046\,
            in1 => \N__40384\,
            in2 => \N__42009\,
            in3 => \N__40365\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49892\,
            ce => 'H',
            sr => \N__49475\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__40382\,
            in1 => \N__42555\,
            in2 => \N__40366\,
            in3 => \N__42484\,
            lcout => \phase_controller_inst2.start_timer_tr_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__40330\,
            in1 => \N__43307\,
            in2 => \N__42252\,
            in3 => \N__40306\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44899\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40288\,
            in2 => \_gnd_net_\,
            in3 => \N__40273\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40270\,
            in2 => \_gnd_net_\,
            in3 => \N__40255\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40252\,
            in2 => \_gnd_net_\,
            in3 => \N__40240\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42856\,
            in2 => \_gnd_net_\,
            in3 => \N__40237\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40465\,
            in2 => \N__42811\,
            in3 => \N__40234\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42760\,
            in2 => \N__40497\,
            in3 => \N__40792\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40469\,
            in2 => \N__42718\,
            in3 => \N__40399\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42670\,
            in2 => \_gnd_net_\,
            in3 => \N__40387\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42625\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42583\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43132\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43084\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43036\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43003\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42976\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42949\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_28_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42922\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43369\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43276\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40804\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48320\,
            in1 => \N__43743\,
            in2 => \_gnd_net_\,
            in3 => \N__43722\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43207\,
            in1 => \N__43605\,
            in2 => \_gnd_net_\,
            in3 => \N__48156\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45450\,
            in1 => \N__43414\,
            in2 => \N__45943\,
            in3 => \N__43472\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45513\,
            in1 => \N__45578\,
            in2 => \N__43895\,
            in3 => \N__48421\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40903\,
            in1 => \N__40897\,
            in2 => \N__40891\,
            in3 => \N__40888\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43507\,
            in1 => \N__48155\,
            in2 => \_gnd_net_\,
            in3 => \N__43481\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__46181\,
            in1 => \N__41444\,
            in2 => \_gnd_net_\,
            in3 => \N__40882\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__40833\,
            in1 => \N__45871\,
            in2 => \N__40861\,
            in3 => \N__45855\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__45870\,
            in1 => \N__40860\,
            in2 => \N__45859\,
            in3 => \N__40834\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45471\,
            in1 => \N__45446\,
            in2 => \_gnd_net_\,
            in3 => \N__48153\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48154\,
            in1 => \N__43189\,
            in2 => \_gnd_net_\,
            in3 => \N__43572\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47296\,
            in1 => \N__47334\,
            in2 => \_gnd_net_\,
            in3 => \N__48173\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__45825\,
            sr => \N__49381\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__43913\,
            in1 => \_gnd_net_\,
            in2 => \N__43896\,
            in3 => \N__48175\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__45825\,
            sr => \N__49381\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44188\,
            in1 => \N__44223\,
            in2 => \_gnd_net_\,
            in3 => \N__48171\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__45825\,
            sr => \N__49381\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43488\,
            in1 => \N__43505\,
            in2 => \_gnd_net_\,
            in3 => \N__48174\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__45825\,
            sr => \N__49381\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44167\,
            in1 => \N__44131\,
            in2 => \_gnd_net_\,
            in3 => \N__48172\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49993\,
            ce => \N__45825\,
            sr => \N__49381\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__41031\,
            in1 => \N__41008\,
            in2 => \N__41059\,
            in3 => \N__41068\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41067\,
            in1 => \N__41058\,
            in2 => \N__41035\,
            in3 => \N__41007\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48328\,
            in1 => \N__43453\,
            in2 => \_gnd_net_\,
            in3 => \N__43422\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49981\,
            ce => \N__45823\,
            sr => \N__49388\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__40969\,
            in1 => \N__40944\,
            in2 => \N__40924\,
            in3 => \N__41353\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41352\,
            in1 => \N__40968\,
            in2 => \N__40948\,
            in3 => \N__40920\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48267\,
            in1 => \N__47189\,
            in2 => \_gnd_net_\,
            in3 => \N__47154\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47190\,
            in1 => \_gnd_net_\,
            in2 => \N__41362\,
            in3 => \N__48269\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49971\,
            ce => \N__45797\,
            sr => \N__49395\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48268\,
            in1 => \N__45613\,
            in2 => \_gnd_net_\,
            in3 => \N__45582\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49971\,
            ce => \N__45797\,
            sr => \N__49395\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48318\,
            in1 => \N__41445\,
            in2 => \_gnd_net_\,
            in3 => \N__41405\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41516\,
            in1 => \N__41493\,
            in2 => \_gnd_net_\,
            in3 => \N__48317\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41802\,
            in2 => \_gnd_net_\,
            in3 => \N__41834\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__41765\,
            in1 => \_gnd_net_\,
            in2 => \N__41344\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41766\,
            in2 => \_gnd_net_\,
            in3 => \N__41328\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41308\,
            in2 => \_gnd_net_\,
            in3 => \N__42146\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__41587\,
            in1 => \N__41557\,
            in2 => \N__41542\,
            in3 => \N__41537\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49407\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__46975\,
            in1 => \N__47014\,
            in2 => \N__46030\,
            in3 => \N__46865\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49407\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__46549\,
            in1 => \N__46569\,
            in2 => \N__41383\,
            in3 => \N__41455\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41454\,
            in1 => \N__46548\,
            in2 => \N__46573\,
            in3 => \N__41379\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41517\,
            in1 => \N__41494\,
            in2 => \_gnd_net_\,
            in3 => \N__48389\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__47916\,
            sr => \N__49414\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48385\,
            in1 => \N__41446\,
            in2 => \_gnd_net_\,
            in3 => \N__41406\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__47916\,
            sr => \N__49414\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46147\,
            in1 => \N__48390\,
            in2 => \_gnd_net_\,
            in3 => \N__46185\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__47916\,
            sr => \N__49414\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41370\,
            in1 => \N__46498\,
            in2 => \N__46528\,
            in3 => \N__41850\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__46524\,
            in1 => \N__46497\,
            in2 => \N__41854\,
            in3 => \N__41371\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41902\,
            in2 => \N__48400\,
            in3 => \N__41884\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__47916\,
            sr => \N__49414\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42093\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49420\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__41646\,
            in1 => \N__41761\,
            in2 => \N__41803\,
            in3 => \N__41841\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49420\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41794\,
            in2 => \_gnd_net_\,
            in3 => \N__42086\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__41814\,
            in1 => \N__41793\,
            in2 => \_gnd_net_\,
            in3 => \N__42085\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41642\,
            in2 => \_gnd_net_\,
            in3 => \N__41598\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__41619\,
            in1 => \N__41734\,
            in2 => \_gnd_net_\,
            in3 => \N__41680\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.state_3_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__42435\,
            in1 => \N__41719\,
            in2 => \N__42118\,
            in3 => \N__44683\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.state_0_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__41679\,
            in1 => \N__41599\,
            in2 => \N__41650\,
            in3 => \N__41618\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst2.start_timer_hc_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__44733\,
            in1 => \N__42523\,
            in2 => \N__42067\,
            in3 => \N__42140\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.start_timer_tr_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__42111\,
            in1 => \N__42100\,
            in2 => \N__42094\,
            in3 => \N__44734\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42033\,
            in2 => \_gnd_net_\,
            in3 => \N__41989\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__42554\,
            in1 => \N__44671\,
            in2 => \N__42501\,
            in3 => \N__44659\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49454\
        );

    \phase_controller_inst1.state_4_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44795\,
            in2 => \_gnd_net_\,
            in3 => \N__44729\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49454\
        );

    \phase_controller_inst2.start_timer_tr_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__44728\,
            in1 => \N__42058\,
            in2 => \N__46939\,
            in3 => \N__44638\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49454\
        );

    \phase_controller_inst2.state_3_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__42045\,
            in1 => \N__44682\,
            in2 => \N__42005\,
            in3 => \N__44637\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49454\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41971\,
            in1 => \N__41953\,
            in2 => \N__41938\,
            in3 => \N__41920\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42577\,
            in1 => \N__42571\,
            in2 => \N__42565\,
            in3 => \N__42562\,
            lcout => \current_shift_inst.PI_CTRL.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__42556\,
            in1 => \N__42491\,
            in2 => \_gnd_net_\,
            in3 => \N__42516\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49893\,
            ce => 'H',
            sr => \N__49476\
        );

    \phase_controller_inst1.test22_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__42387\,
            in1 => \N__42436\,
            in2 => \N__44740\,
            in3 => \N__44804\,
            lcout => test22_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49893\,
            ce => 'H',
            sr => \N__49476\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50241\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => 'H',
            sr => \N__49486\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42192\,
            in2 => \_gnd_net_\,
            in3 => \N__44844\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__45268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42180\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__42181\,
            in1 => \N__45256\,
            in2 => \N__42172\,
            in3 => \N__44971\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45300\,
            in2 => \_gnd_net_\,
            in3 => \N__42159\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__45200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43242\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42909\,
            in2 => \_gnd_net_\,
            in3 => \N__45336\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42898\,
            in2 => \N__42877\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_16_27_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42850\,
            in2 => \N__42832\,
            in3 => \N__42802\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42799\,
            in2 => \N__42781\,
            in3 => \N__42754\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42751\,
            in2 => \N__42733\,
            in3 => \N__42709\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42706\,
            in2 => \N__42691\,
            in3 => \N__42664\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42661\,
            in2 => \N__42643\,
            in3 => \N__42619\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42616\,
            in2 => \N__42604\,
            in3 => \N__43171\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43168\,
            in2 => \N__43153\,
            in3 => \N__43126\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43123\,
            in2 => \N__43108\,
            in3 => \N__43078\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_16_28_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43075\,
            in2 => \N__43057\,
            in3 => \N__43030\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43327\,
            in2 => \N__43027\,
            in3 => \N__42997\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42994\,
            in2 => \N__43340\,
            in3 => \N__42970\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43331\,
            in2 => \N__42967\,
            in3 => \N__42943\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42940\,
            in2 => \N__43341\,
            in3 => \N__42916\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43335\,
            in2 => \N__43390\,
            in3 => \N__43363\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43360\,
            in2 => \N__43342\,
            in3 => \N__43270\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43267\,
            in1 => \N__43261\,
            in2 => \_gnd_net_\,
            in3 => \N__43249\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_16_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__43246\,
            in1 => \N__45201\,
            in2 => \N__44972\,
            in3 => \N__45178\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_16_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__44945\,
            in1 => \N__45130\,
            in2 => \N__45154\,
            in3 => \N__45247\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43206\,
            in1 => \N__43606\,
            in2 => \_gnd_net_\,
            in3 => \N__48170\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__47911\,
            sr => \N__49374\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43188\,
            in1 => \N__43573\,
            in2 => \_gnd_net_\,
            in3 => \N__48169\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50015\,
            ce => \N__47911\,
            sr => \N__49374\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43821\,
            in1 => \N__43858\,
            in2 => \_gnd_net_\,
            in3 => \N__48221\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48223\,
            in1 => \N__43915\,
            in2 => \_gnd_net_\,
            in3 => \N__43888\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43990\,
            in2 => \_gnd_net_\,
            in3 => \N__44065\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48222\,
            in1 => \N__43689\,
            in2 => \_gnd_net_\,
            in3 => \N__43662\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43598\,
            in1 => \N__43565\,
            in2 => \N__44137\,
            in3 => \N__44215\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__45398\,
            in1 => \N__43772\,
            in2 => \N__43534\,
            in3 => \N__43531\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__47543\,
            in1 => \N__43525\,
            in2 => \N__43519\,
            in3 => \N__43516\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44216\,
            in1 => \_gnd_net_\,
            in2 => \N__43510\,
            in3 => \N__44186\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48157\,
            in1 => \N__43506\,
            in2 => \_gnd_net_\,
            in3 => \N__43489\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45900\,
            in1 => \N__45941\,
            in2 => \_gnd_net_\,
            in3 => \N__48163\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48159\,
            in1 => \N__43449\,
            in2 => \_gnd_net_\,
            in3 => \N__43426\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47292\,
            in1 => \N__47335\,
            in2 => \_gnd_net_\,
            in3 => \N__48162\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__48158\,
            in1 => \N__43914\,
            in2 => \N__43897\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43857\,
            in1 => \N__43817\,
            in2 => \_gnd_net_\,
            in3 => \N__48160\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43800\,
            in1 => \N__48164\,
            in2 => \_gnd_net_\,
            in3 => \N__43780\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43744\,
            in1 => \N__43721\,
            in2 => \_gnd_net_\,
            in3 => \N__48161\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50004\,
            ce => \N__47912\,
            sr => \N__49379\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__46626\,
            in1 => \N__46605\,
            in2 => \N__43618\,
            in3 => \N__43627\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__43626\,
            in1 => \N__46627\,
            in2 => \N__46606\,
            in3 => \N__43614\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48270\,
            in1 => \N__43685\,
            in2 => \_gnd_net_\,
            in3 => \N__43663\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49994\,
            ce => \N__47913\,
            sr => \N__49382\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47362\,
            in1 => \N__47397\,
            in2 => \_gnd_net_\,
            in3 => \N__48273\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49994\,
            ce => \N__47913\,
            sr => \N__49382\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44224\,
            in1 => \N__44187\,
            in2 => \_gnd_net_\,
            in3 => \N__48271\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49994\,
            ce => \N__47913\,
            sr => \N__49382\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44163\,
            in1 => \N__44136\,
            in2 => \_gnd_net_\,
            in3 => \N__48272\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49994\,
            ce => \N__47913\,
            sr => \N__49382\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__46098\,
            in1 => \N__46336\,
            in2 => \N__46363\,
            in3 => \N__46114\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44098\,
            in1 => \N__44071\,
            in2 => \_gnd_net_\,
            in3 => \N__48275\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49982\,
            ce => \N__47915\,
            sr => \N__49389\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44034\,
            in1 => \N__48274\,
            in2 => \_gnd_net_\,
            in3 => \N__44002\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49982\,
            ce => \N__47915\,
            sr => \N__49389\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46016\,
            in1 => \N__43945\,
            in2 => \N__43960\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43927\,
            in2 => \N__43939\,
            in3 => \N__46002\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43921\,
            in2 => \N__45415\,
            in3 => \N__45972\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45957\,
            in1 => \N__44371\,
            in2 => \N__44359\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45349\,
            in2 => \N__44347\,
            in3 => \N__46311\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46297\,
            in1 => \N__44338\,
            in2 => \N__44329\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44320\,
            in2 => \N__44314\,
            in3 => \N__46278\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44305\,
            in2 => \N__44299\,
            in3 => \N__46264\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44287\,
            in2 => \N__44278\,
            in3 => \N__46245\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44269\,
            in2 => \N__44260\,
            in3 => \N__46230\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46215\,
            in1 => \N__44248\,
            in2 => \N__44236\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46200\,
            in1 => \N__44452\,
            in2 => \N__44464\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44434\,
            in2 => \N__44446\,
            in3 => \N__46473\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46458\,
            in1 => \N__47143\,
            in2 => \N__44428\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46443\,
            in1 => \N__44419\,
            in2 => \N__44410\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47206\,
            in2 => \N__47059\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46042\,
            in2 => \N__45628\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44401\,
            in2 => \N__46081\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44392\,
            in2 => \N__44383\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47734\,
            in2 => \N__47794\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44524\,
            in2 => \N__44518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44509\,
            in2 => \N__44503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47470\,
            in2 => \N__47410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44494\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46902\,
            in2 => \_gnd_net_\,
            in3 => \N__47030\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44491\,
            in3 => \N__46967\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => 'H',
            sr => \N__49421\
        );

    \phase_controller_inst1.test_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__44475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44735\,
            lcout => test_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => 'H',
            sr => \N__49429\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__44657\,
            in1 => \N__46968\,
            in2 => \N__46911\,
            in3 => \N__47035\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => 'H',
            sr => \N__49429\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44777\,
            in2 => \_gnd_net_\,
            in3 => \N__44713\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44670\,
            in2 => \_gnd_net_\,
            in3 => \N__44658\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44611\,
            in2 => \_gnd_net_\,
            in3 => \N__44629\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44587\,
            in2 => \_gnd_net_\,
            in3 => \N__44605\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44566\,
            in2 => \_gnd_net_\,
            in3 => \N__44581\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44548\,
            in2 => \_gnd_net_\,
            in3 => \N__44560\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44530\,
            in2 => \_gnd_net_\,
            in3 => \N__44542\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45100\,
            in2 => \_gnd_net_\,
            in3 => \N__45115\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45079\,
            in2 => \_gnd_net_\,
            in3 => \N__45094\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45058\,
            in2 => \_gnd_net_\,
            in3 => \N__45073\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45034\,
            in2 => \_gnd_net_\,
            in3 => \N__45052\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_17_27_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45010\,
            in2 => \_gnd_net_\,
            in3 => \N__45028\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46649\,
            in2 => \_gnd_net_\,
            in3 => \N__44995\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__44949\,
            in1 => \N__44898\,
            in2 => \_gnd_net_\,
            in3 => \N__44854\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44840\,
            in2 => \_gnd_net_\,
            in3 => \N__44815\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45332\,
            in2 => \_gnd_net_\,
            in3 => \N__45307\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45296\,
            in2 => \_gnd_net_\,
            in3 => \N__45271\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45267\,
            in2 => \_gnd_net_\,
            in3 => \N__45250\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_17_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45128\,
            in2 => \_gnd_net_\,
            in3 => \N__45241\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_17_28_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45238\,
            in2 => \_gnd_net_\,
            in3 => \N__45205\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45202\,
            in2 => \_gnd_net_\,
            in3 => \N__45172\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45169\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__45129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45153\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45893\,
            in1 => \N__45942\,
            in2 => \_gnd_net_\,
            in3 => \N__48276\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45605\,
            in1 => \N__45583\,
            in2 => \_gnd_net_\,
            in3 => \N__48152\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47271\,
            in1 => \N__47244\,
            in2 => \_gnd_net_\,
            in3 => \N__48242\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50016\,
            ce => \N__45836\,
            sr => \N__49375\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48459\,
            in1 => \N__48432\,
            in2 => \_gnd_net_\,
            in3 => \N__48243\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50016\,
            ce => \N__45836\,
            sr => \N__49375\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__46065\,
            in1 => \N__46419\,
            in2 => \N__46393\,
            in3 => \N__46053\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45606\,
            in1 => \N__45574\,
            in2 => \_gnd_net_\,
            in3 => \N__48168\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => \N__47914\,
            sr => \N__49377\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48165\,
            in1 => \N__45541\,
            in2 => \_gnd_net_\,
            in3 => \N__45514\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => \N__47914\,
            sr => \N__49377\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48166\,
            in1 => \N__45475\,
            in2 => \_gnd_net_\,
            in3 => \N__45451\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => \N__47914\,
            sr => \N__49377\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48167\,
            in1 => \N__45403\,
            in2 => \_gnd_net_\,
            in3 => \N__45373\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50011\,
            ce => \N__47914\,
            sr => \N__49377\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48277\,
            in1 => \N__46186\,
            in2 => \_gnd_net_\,
            in3 => \N__46136\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__46110\,
            in1 => \N__46335\,
            in2 => \N__46099\,
            in3 => \N__46359\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47270\,
            in1 => \N__47243\,
            in2 => \_gnd_net_\,
            in3 => \N__48278\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__46066\,
            in1 => \N__46392\,
            in2 => \N__46423\,
            in3 => \N__46054\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46029\,
            in2 => \N__46999\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46824\,
            in1 => \N__46003\,
            in2 => \_gnd_net_\,
            in3 => \N__45991\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__46866\,
            in1 => \N__45988\,
            in2 => \N__45976\,
            in3 => \N__45961\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46825\,
            in1 => \N__45958\,
            in2 => \_gnd_net_\,
            in3 => \N__45946\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46867\,
            in1 => \N__46312\,
            in2 => \_gnd_net_\,
            in3 => \N__46300\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46826\,
            in1 => \N__46296\,
            in2 => \_gnd_net_\,
            in3 => \N__46282\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46868\,
            in1 => \N__46279\,
            in2 => \_gnd_net_\,
            in3 => \N__46267\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46827\,
            in1 => \N__46263\,
            in2 => \_gnd_net_\,
            in3 => \N__46249\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49995\,
            ce => 'H',
            sr => \N__49383\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46835\,
            in1 => \N__46246\,
            in2 => \_gnd_net_\,
            in3 => \N__46234\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46820\,
            in1 => \N__46231\,
            in2 => \_gnd_net_\,
            in3 => \N__46219\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46832\,
            in1 => \N__46216\,
            in2 => \_gnd_net_\,
            in3 => \N__46204\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46821\,
            in1 => \N__46201\,
            in2 => \_gnd_net_\,
            in3 => \N__46189\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46833\,
            in1 => \N__46474\,
            in2 => \_gnd_net_\,
            in3 => \N__46462\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46822\,
            in1 => \N__46459\,
            in2 => \_gnd_net_\,
            in3 => \N__46447\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46834\,
            in1 => \N__46444\,
            in2 => \_gnd_net_\,
            in3 => \N__46432\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46823\,
            in1 => \N__47078\,
            in2 => \_gnd_net_\,
            in3 => \N__46429\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49983\,
            ce => 'H',
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46828\,
            in1 => \N__47126\,
            in2 => \_gnd_net_\,
            in3 => \N__46426\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46869\,
            in1 => \N__46418\,
            in2 => \_gnd_net_\,
            in3 => \N__46396\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46829\,
            in1 => \N__46388\,
            in2 => \_gnd_net_\,
            in3 => \N__46366\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46870\,
            in1 => \N__46358\,
            in2 => \_gnd_net_\,
            in3 => \N__46339\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46830\,
            in1 => \N__46334\,
            in2 => \_gnd_net_\,
            in3 => \N__46315\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46871\,
            in1 => \N__46625\,
            in2 => \_gnd_net_\,
            in3 => \N__46609\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46831\,
            in1 => \N__46596\,
            in2 => \_gnd_net_\,
            in3 => \N__46582\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46872\,
            in1 => \N__47769\,
            in2 => \_gnd_net_\,
            in3 => \N__46579\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49972\,
            ce => 'H',
            sr => \N__49396\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46842\,
            in1 => \N__47754\,
            in2 => \_gnd_net_\,
            in3 => \N__46576\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46836\,
            in1 => \N__46568\,
            in2 => \_gnd_net_\,
            in3 => \N__46552\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46843\,
            in1 => \N__46547\,
            in2 => \_gnd_net_\,
            in3 => \N__46531\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46837\,
            in1 => \N__46523\,
            in2 => \_gnd_net_\,
            in3 => \N__46501\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46844\,
            in1 => \N__46496\,
            in2 => \_gnd_net_\,
            in3 => \N__46477\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46838\,
            in1 => \N__47447\,
            in2 => \_gnd_net_\,
            in3 => \N__47041\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46845\,
            in1 => \N__47426\,
            in2 => \_gnd_net_\,
            in3 => \N__47038\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49401\
        );

    \phase_controller_inst2.stoper_tr.running_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__46987\,
            in1 => \N__46966\,
            in2 => \N__46912\,
            in3 => \N__47034\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => 'H',
            sr => \N__49408\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46965\,
            in2 => \_gnd_net_\,
            in3 => \N__47010\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__46903\,
            in1 => \N__46986\,
            in2 => \_gnd_net_\,
            in3 => \N__46940\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46941\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46904\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46726\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49422\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46674\,
            in2 => \_gnd_net_\,
            in3 => \N__46653\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50023\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47357\,
            in1 => \N__47398\,
            in2 => \_gnd_net_\,
            in3 => \N__48315\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47291\,
            in1 => \N__47333\,
            in2 => \_gnd_net_\,
            in3 => \N__48297\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48298\,
            in1 => \N__47272\,
            in2 => \_gnd_net_\,
            in3 => \N__47248\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50017\,
            ce => \N__47917\,
            sr => \N__49380\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__47932\,
            in1 => \N__47103\,
            in2 => \N__47131\,
            in3 => \N__47088\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48299\,
            in1 => \N__47194\,
            in2 => \_gnd_net_\,
            in3 => \N__47158\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50012\,
            ce => \N__47918\,
            sr => \N__49384\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47492\,
            in1 => \N__47544\,
            in2 => \_gnd_net_\,
            in3 => \N__48282\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__47127\,
            in1 => \N__47104\,
            in2 => \N__47089\,
            in3 => \N__47931\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48283\,
            in1 => \N__47624\,
            in2 => \_gnd_net_\,
            in3 => \N__47601\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48647\,
            in1 => \N__48624\,
            in2 => \_gnd_net_\,
            in3 => \N__48284\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47715\,
            in1 => \N__47694\,
            in2 => \_gnd_net_\,
            in3 => \N__48353\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__47554\,
            in1 => \N__47641\,
            in2 => \N__47779\,
            in3 => \N__47753\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__47640\,
            in1 => \N__47775\,
            in2 => \N__47755\,
            in3 => \N__47553\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48354\,
            in1 => \N__47711\,
            in2 => \_gnd_net_\,
            in3 => \N__47695\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__47920\,
            sr => \N__49402\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47625\,
            in1 => \N__47602\,
            in2 => \_gnd_net_\,
            in3 => \N__48356\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__47920\,
            sr => \N__49402\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48355\,
            in1 => \N__47545\,
            in2 => \_gnd_net_\,
            in3 => \N__47496\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__47920\,
            sr => \N__49402\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__48579\,
            in1 => \N__47451\,
            in2 => \N__47431\,
            in3 => \N__47460\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__47461\,
            in1 => \N__48580\,
            in2 => \N__47452\,
            in3 => \N__47430\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48648\,
            in1 => \N__48625\,
            in2 => \_gnd_net_\,
            in3 => \N__48357\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49984\,
            ce => \N__47920\,
            sr => \N__49402\
        );

    \delay_measurement_inst.stop_timer_tr_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48494\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__49437\
        );

    \delay_measurement_inst.start_timer_tr_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48493\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__49437\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48458\,
            in1 => \N__48431\,
            in2 => \_gnd_net_\,
            in3 => \N__48316\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48460\,
            in1 => \N__48436\,
            in2 => \_gnd_net_\,
            in3 => \N__48352\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50018\,
            ce => \N__47919\,
            sr => \N__49391\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47884\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47860\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49482\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__48667\,
            in1 => \N__48721\,
            in2 => \N__48880\,
            in3 => \N__48661\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48897\,
            in2 => \_gnd_net_\,
            in3 => \N__48773\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50405\,
            in2 => \_gnd_net_\,
            in3 => \N__50297\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__50345\,
            in1 => \N__50505\,
            in2 => \N__48691\,
            in3 => \N__50178\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__50243\,
            in1 => \N__48683\,
            in2 => \N__48923\,
            in3 => \N__50123\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__50242\,
            in1 => \N__48684\,
            in2 => \_gnd_net_\,
            in3 => \N__50122\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__50244\,
            in1 => \N__48688\,
            in2 => \N__48924\,
            in3 => \N__50124\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50468\,
            in2 => \_gnd_net_\,
            in3 => \N__50264\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__50321\,
            in1 => \N__50375\,
            in2 => \N__48670\,
            in3 => \N__50039\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__50430\,
            in1 => \N__48954\,
            in2 => \_gnd_net_\,
            in3 => \N__48819\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50322\,
            in1 => \N__50376\,
            in2 => \N__50473\,
            in3 => \N__50040\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__48655\,
            in1 => \N__48720\,
            in2 => \N__48876\,
            in3 => \N__50265\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__50174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50412\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50298\,
            in1 => \N__50352\,
            in2 => \N__48997\,
            in3 => \N__50501\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__50240\,
            in1 => \N__48994\,
            in2 => \N__48988\,
            in3 => \N__50063\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__48786\,
            in1 => \N__48798\,
            in2 => \N__48985\,
            in3 => \N__48774\,
            lcout => \current_shift_inst.PI_CTRL.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48976\,
            in2 => \_gnd_net_\,
            in3 => \N__50443\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__48940\,
            in1 => \N__48931\,
            in2 => \N__48925\,
            in3 => \N__50079\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48841\,
            in2 => \_gnd_net_\,
            in3 => \N__50442\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__48805\,
            in1 => \N__48787\,
            in2 => \_gnd_net_\,
            in3 => \N__48775\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__50245\,
            in1 => \N__50121\,
            in2 => \N__50506\,
            in3 => \N__50078\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50452\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50441\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49490\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010100"
        )
    port map (
            in0 => \N__50239\,
            in1 => \N__50416\,
            in2 => \N__50143\,
            in3 => \N__50083\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49494\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110110000"
        )
    port map (
            in0 => \N__50082\,
            in1 => \N__50238\,
            in2 => \N__50359\,
            in3 => \N__50141\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49494\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110110000"
        )
    port map (
            in0 => \N__50080\,
            in1 => \N__50236\,
            in2 => \N__50305\,
            in3 => \N__50140\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49494\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010100"
        )
    port map (
            in0 => \N__50237\,
            in1 => \N__50179\,
            in2 => \N__50142\,
            in3 => \N__50081\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49494\
        );
end \INTERFACE\;
